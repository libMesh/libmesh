netcdf test_one_var {
variables:
  int t;
data:
  t = 17;
}
