netcdf tst_special_atts {
types:
  compound obs_t {
    byte day ;
    short elev ;
    int count ;
    float relhum ;
    double time ;
    ubyte category ;
    ushort id ;
    uint particularity ;
    int64 attention_span ;
  }; // obs_t
dimensions:
	dim1 = 10 ;
	dim2 = 20 ;
	dim3 = 30 ;
variables:
	int var1(dim1) ;
		var1:_Storage = "contiguous" ;
		var1:_Endianness = "little" ;
	int var2(dim1, dim2) ;
		var2:_Storage = "chunked" ;
		var2:_ChunkSizes = 6, 7 ;
		var2:_Fletcher32 = "true" ;
		var2:_Endianness = "big" ;
	int var3(dim1, dim2, dim3) ;
		var3:_Storage = "chunked" ;
		var3:_ChunkSizes = 6, 7, 8 ;
		var3:_DeflateLevel = 2 ;
		var3:_Endianness = "little" ;
	int var4(dim1, dim2, dim3) ;
		var4:_Storage = "chunked" ;
		var4:_ChunkSizes = 6, 7, 8 ;
		var4:_DeflateLevel = 2 ;
		var4:_Shuffle = "true" ;
		var4:_Endianness = "little" ;
		var4:_NoFill = "true" ;
	obs_t var5(dim1) ;
		var5:_Storage = "chunked" ;
		var5:_ChunkSizes = 6 ;
		var5:_DeflateLevel = 2 ;
		var5:_Shuffle = "true" ;
		var5:_Fletcher32 = "true" ;
		var5:_NoFill = "true" ;

// global attributes:
 		:_NCProperties = "version=2,netcdf=4.6.2-development,hdf5=1.10.1" ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
data:
}
