netcdf ref_typescope {

group: f {
types:
  opaque(3) op_t1;
} // group f

group: g {
  types:
    opaque(4) op_t2 ;
  variables:
      op_t1 v1 ; // use /f/op_t1
  data:

   v1 = 0X000000  ;

  group: h {
    types:
      opaque(4) op_t3 ;
    variables:
      op_t2 v2 ; // use /g/op_t2
    data:

     v2 = 0X00000000 ;
  } // group h

  group: i {
    types:
      opaque(4) op_t2 ;
    variables:
      op_t3 v2 ; // use /g/h/op_t3
    data:

     v2 = 0X00000000 ;
  } // group i
} // group g

group: j {
  variables:
    op_t3 v2 ; // use /g/h/op_t3
  data:

   v2 = 0X00000000 ;
} // group j
}
