netcdf test_vlen3 {

types:
  int(*) v_t;
  compound c_t {v_t f1;};

variables:
  c_t v1;  

data:
  v1 = {{1, 3, 5, 7}} ;
}

