netcdf test_vlen5 {

types:
  int(*) v_t;
  compound c_t {v_t v;};

dimensions:
  d2=2;

variables:
  c_t v1(d2);  

data:
  v1 = {{1, 3, 5, 7}},{{100,200}} ;
}

