netcdf tst_chunks {
dimensions:
	dim1 = 32 ;
	dim2 = 90 ;
	dim3 = 91 ;
variables:
	float var_contiguous(dim1, dim2, dim3) ;
		var_contiguous:_Storage = "contiguous" ;
		var_contiguous:_Endianness = "little" ;
	float var_chunked(dim1, dim2, dim3) ;
		var_chunked:_Storage = "chunked" ;
		var_chunked:_ChunkSizes = 8, 10, 13 ;
		var_chunked:_Endianness = "little" ;
	float var_compressed(dim1, dim2, dim3) ;
		var_compressed:_Storage = "chunked" ;
		var_compressed:_ChunkSizes = 8, 10, 13 ;
		var_compressed:_DeflateLevel = 1 ;
		var_compressed:_Endianness = "little" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.2-development|hdf5libversion=1.8.17" ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4 classic model" ;
}
