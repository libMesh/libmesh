netcdf tst_long_charconst {
dimensions:
	obs = 60000 ;
variables:
	char PRCP_MFLAG(obs) ;
data:

 PRCP_MFLAG = " PPPP PP PP PP PPP PPPPPPPPP PP P PPP PPP P P PP PPP PPPPP                               PPPPPPP  P P P PPPPP  PPPP P P PP P PPPPPP PP TTPPPP PPPPP PP   T                          P  PPP  PPPPP P P PPPPPPP PPPP PPPP  PPPPP PPPP PP PPP PPPP PPP PPPPPPPPPPPP  PPPPPP P P PPP                                                             PP  PPPP PPPP  PPPPP PPPPP PP PPPP P PPP PPPP PP P PPP P PP PPPP PPPPP PP P PP PPP PPP PPPPPPPP PPP PPPP PP P P PP PP PP                              PPPPP PPPPPPPPP PPPP P PPPPP P PPP PPPPPPP  P PP P PPPPP PPPPPPPPPPP P PPPPPPP P PPPPPPPPP PPPP  PPPP PP PPPPPPPPPPP PP PP PP P PPP PPPP PPP PP P PPPPPPPP PPPPPP PP PPPPPPPPPPPPPP PPPPPPPPPP PP P PPP PPPP PPPP PP PPP PPPP PPPPP PPPPPPPPPPPPPP P PPPPPP PPP PP PPPPPPPPPPPPPPPPP PPPP PPPP PPPPPPPPPPPPPPPP PP PP  PPPP P P P PPP PPP  PPPP         T                     PPPP PPPPPPPP PPPPPPPPPPP PPPPPPPPP  PPPPPPPP PPPPPPPPPPPPPP PPPPPP  PPPPPPPPP PPPPPP PPPPP                               P PPPPPPP PPPP P PP PPPP  PPPP PPPPPP PPPPPPPPPPP PPPP PPPP PPPPPPPPPPPPPPPPPPPP PPP  PPPPP  PPPP  P PPPP PPPP PPPPPPPPP PPPPPP PPPP PPP PP PPP PPPPPP PP PPP PPP PPPPPPPP PPPP PPPPPPPP P PPPPPP PPPPP PP PPP PP PPPPPPPPPP   PPP PP P P PPP PP PPP PPPPPPPPPPP PPPPPPP   PPPPPPPPP P PPPPPPPPP PPP PPPPPPPPPP PPP PPPPPPPP PPPPPPPPP PPPPPPPPPPPP PPPPPP PPPPPPPPP PPPPPPP PPPPPPPP PPPPPP PPPPPPPPPP PPPPPPPPP PPP  PPP PPPP P PP PPPPP                             PTTP PTPPP PPP PPP PPPP   P PPP PPPPP PP   P P PPPPPP   PPPPPPPPPPPPPPP PP PPPP PP PPPPP PP                                                                                           PPPPP PPP PPP PP   PP   P PPP PPP PPPPPPP PPPP PP P PPPPPPPPPP  PPP  TPPPPPPPPPPPPPPPPP  PP  PPPP PPP PP PPPP  PP  P PPPPP P  PPPP  PPPPP  PP P P PPPP  P   PPPPPPPP PPPPPPPP PPPP    PPPP PPPPPPPP PPPPPPPPP PPPPPP P PP P PP PPPPPPPPP    PPPPPPPP PPPPPPPPPP PPP PP   PPPPPPPPPPPPPP  PP  PPPPP   P PPPPPP PPP PPP PPP PPP      PPPPPPTPT PP P PP  PPPPPPPPPPPPPPTPP PPPPPP PPP PPP PP  PPPP PPPPPPPPPPP PPPPPP P TPTTPPPPP PPP PP PPPP PP P  P P PPPP PP  PPPPP  PPPTP PP PP PP PP PPPP PPPPP PPP PP PPPP PPP  PPPPP PPPPPP PPP PPPP P PPP  PPTPPP PP PPP PPPPPPP        T                     PPP PPP PPPPPPPPPPP PPPPPP  PPPPPPPP  PP P PPPPP  P    P PPPP P  PPPP  PPP PPTPPPPP PPPPPP PPPP PP PPPP PPPPPPPPPP  P PPTPP PPP  PPPPPP T TPP TPPTPP PPP PPPP PP PPPPP TPPPPPP PPPP  P P  P PP P PPPP  P  PPPPP P  T        T                      PPPPPPPPPPTPPP PPPPTPPPPPPPPPPPP  PPPPPPPTP PPPPPPT      PPP PPPP   P P PPPTT P PPTPP   PPPPTPPPP PPPPPPPPPPPPPPPPPPPPP PPPPPPPPPPT PPPPPPPPPPPPPPT T  PPPPPPPPPPPPPPP PPPTPPPPPPPPPPPPPPPTPP PPP PPPPP TPPP PP PPPPPPPPPP P PPPPPP PT PPPPP PPPPP PTPPPPPT  T PP PP PP PTPP PPPPPP  PTPPP PP PPPPP PPPPT PP PPPPTPPPPPP PPPP PPPPP  P PPP PPT PPPPPTPP PPPPPPPPPPP PPPT PPPPPP  PPP    P   P PPPPPPPPPP PPP PPP PPPPPPP PPPPPPPT PPPPPPPPTPP PP PPPPPTPP PPPPPPPPPPPPPPPPPPPPPPPP PPPPP PPPPPPP PP PPPPPPPPPPPPP PP PPPTPP P TPPPTPPPP PPPPPP PPPPPPP PPPPPT  PPPPPPPTPPP PPPPP PPTPPPPPPPP PTP PPPPPPP PPPPPPP PPP PP PPP PP  P PP PPPPPTP PPPPP PPTP PPPPTPP PPPPTPP  PPPPPPPPTPPPPPPPPPPPPPT P PP PPTPPPP   T PP  PPP PPP PPPP     PPPPP P  P   PPP  PTP P P P T   T     PPPPPPP PPPPP PPP PP P PPPP  PPPPPPPPTPP PPTP PPPTP PPPP  PP PPTPPP P PPP   PP PPPPPPPPPPPPPPPPPPPPPPPPPPPPPP  PPPPPPPPPP  P PP PP PPPPPP  PPPPPPPPPPPPPPPPPPP PPP PTTPT  PPPP TPPPPP PPPPT PPPTP P   TPPPP PP  P PPPPPT PPP P  PPTTP P P  PPPP TPTPP PPPPPPPPPPPTP P PPPP   PPP PPPPPPP P TPPPT  PTT PPPP  PPP  T PPPPPPPPPPPPPPP PPP PPPPP PPPPPPPPPPPP PPPP PPPPPP  P  T PPPPP PP PPPPPPPPPPPPPP P PP PPPPPP P PPPPPPP T PPPPP P P P  PPPPP    P   PP PPPPP P TPP TPPPPT PPPPPP P  PPPP PPP PPP PP     PPPPPPPPPTPPPP PP TP PP PP PPPPP PPP PP              T                PP PPP  PPP PP PPP PPPPPP PP PPPTP PPPPPPPTPPTPPTPP PPPP PPP PP P PP PP PP PPPPP PT  PPP PPP PPPP PPPPP PPT  PPP PPPP P TPPPP    PPP PP   PPPPPPPPPPPTPPPP PP PPPPPPPP  PP PPPPP P P PPPPPPPPPP  PP PP  PP PP PPPPPPPPP PPPPPPTPP PPPP  PPPPPPP PPPTPTPPPP  PPTPPPPP P  PP   PTPPPPPPPPPPPPPPPP PPPPPPPP  PPPPPPP PPPPP PPPPPP PPPPPPPPPPPPP PPP PP PPPPP PPPPPP  PPPP PP PP PPP PPP  PP  PPP P PP P  PP PPPTPP  P PPPP PPPPP PPPTTPPPP PPPPPPPPPP PP   TPPP  PPPP  PP  PPPPPTPPPP      PPTPPP PPP P PPPPPPPTPPTPPT T  PPP    PPP P  PPP PP PPPPPPPPPPPP     PT  PPP PPTPPP PP PPPPP PPPPP PPPPPPP PPPPP PP PT PPPPTPPP PPPP PP PP P PT  PPPP PPPP    PPPPPPPTP   PPP  TPP PPPPPT  PPP   P PPPPPPPPPP  PPPPT  PPPPPPPPPPT PPTTPPPP PPTPPPPPPPPPPTP P TPPPPPPP T PPPPPPTTPPPPPPPPPP PPPPPT PPPPP  PPPTP  P PP TPP PPPPPT PPT PPPP PPPPPP P P PPP P P P                            TTPPPP PP  PPP PPPPPPPPPPPPP PPPPTPP PPP PPPPP  PPP PP P  P  PP PPP P PTP T TPPPPPPPPP  PP PPPPPT PPPPPP  PPPPPPPP PP   P  PPPPPTPPPPPPP PPPPPPPPPPPP PPPPPPPPP PPPPPPPPP   PPPPPPPPTPPPPPP PPPPPP PPPPP  PPTPPPPPPPPPPPP TP    PPP   PPPP P PP PPPP  PPPPPPP PPPP  PPP     P   PPPPP    PP PPPPPPPPP PPPPPPP  PPPPPPPP  PPPPPPPPPPP PPPPPPPPPPPP T                    T    T                          T         T            T   T         T      T      T            T                   T   T               T                   T                                             P T       T T              T                   T   T   T     T        T                        T            T                  T                                                               P                                         TPPPT  T PPPP   P   PPTPPPPP P   TPPPPPPPP  PPPPPPPPPP  PPPPPP  PPP PPP P    T PPPPP  TPPTPPP     PPPPP   PPPPPPPPPP P PPT PPPPP     P   PP P TPPP PPPP TP PTPPPP  PPPPPP  P P     P PPP TPP    PP PT P PPPPPT TT PPP PPPT   PPPP  TP  P  PPPPP  P PPT    PPTPPPP PPT  PT P PP   PP PPPPPP TPPT  TPPPPP  P   PPPPPPP    PT P        PT PPP PPPPPPP TPPP PPP TP TP  TPPPP PPPPPP  TP   PPT P T T     P   PP  PPPPPPP TP  P PPPPPPPPPPPPPTP T  PPPPPPPPPPPPPPPPPTPPPPPPPP PPP                                PP PPPP PPT  TTPPPP  PPP PPPP  PPPP  P   P  PPPPPP PPPPPPPP   PPP PP   PPPPPPPP   PPPP PPT  PP P  PP PPPP PP TP PPPP P       T  T                      T    PPPP   P PPPPPPPP TPP  PPPPPPP  PPP PPPP  PPPPPPP P P  TPPPTPP     P  PPPPPPPPP PP   P   P P PPPP   P  PPPPPPPPPP PPPPTTTP TPP   P PPPPP  PPTT TP PP  PPP PPP PPPPPPP PPPPPPPPPP    PPPPP  P   PP PP  PT P T  PP   TPPPTPP  TPPP PPPP   PTP PPPPP  PP PP  PPPPP  P PPPPPP  PP                            T    P  P   PT P PP  PPPPPP       T   TT             T T     PP    TPPPP PP P  TPPP PPTTPPPP   P   P  P PPPP  P  PPP P   PP    PP PPPPP PPPP  PPPPTP  PPP  PPP P  TP   PPPP PPPPP P  PP   PPTPP PP  PPPPPPPPPPPPPPPPPPPPPPPP    PPPP T PPPPP PPPPPPPPPT PPP PPPPPPP  PPTPPPPPTTTTPPPP P P  P P P  P PPPTPPPPP   PP P  PPP  TPPPT TPPPP  P PPP  PT   P   P T P PPPPPP  TPPP  TT       T            TT       PPPP  P PPPP   PPPPPPPPPPPPPP               TT  T                                                         T    T T       T     T                     T                   T          PPPPPPPPPP PPPTPPPP PP  PPPPTP PPPPP  PPPP PPPPTPPPPP PPP PT PPPP  PPP  PP PPPPP P   PP  P PP  PPPPPPP PPPP  PPTPPPP PPPPP        T    TTT T            PPPPP P P   PPPPPPPP  PPP TP PP  PPP    P PPPPPP   P PP PPPP  PPPPPP  P  PPP PPP  PP      PPP  PPP   PP   PPPP T  PP  PP PP PP PT P PPTPPPTPPPPP PPPPPPPPTP PPPPTP P PPPPPPPPPPP   PPPPPPT P PPP  PPT PP PPP   PPPPP  PPP PPP PPPPPPPPPPPPPPPPPP PPPPPPPPPPPP PT PP PPPPPP P PPPP P                T                                           PT PPPPPP   PP  PPPPPPT P PP PPP  PPPPPP PPP P PPPPPPP  T P               T                  TT   T           T        PPPPPPPP  PPPPPPPPPP P P PPPP PPPP TP   P PP P PPPP  P    PP PPPP PPP PP P PPPPPP PPPPPPPPPPPP PPP  PPPPPPP PPPPPPPPPPPPPPPPP  PPP PPPPP P PPPP    PPPPP P  PP P PPP P   PPPPPPTPTP PPPP     PPPPPPPPP PPPP P PPTPPPPPPPP   PP PPPPPPPP  P  PPTPTPPP         T T T               T PPPP  TP  PPPTP PP P PP PPPP  PP P    P  P PPPTPPPP PP P  PPPPTPPPPPTTPP    PPPPP  PPPPPP  PP    PPPPPPP PPPPPP  PP PPPPPPPPP  PPPPPP   PP  PPPP PPP    PPPPPPPPPPPPT P    P  T PPPPPPP  PPP PP PPPPPPPPPPPPP   P   PPPPP PPPP P  PP  P  P   PPP P TPPPPPPP  PPPP  PP PPPPPP  PP PPTP PTPPPPP  P PPPTP PTPP   PPTP  PTPPTT", "PPP   PPP  PT PPPP  P  T            T    TT  T  T     T                       TT      TP PPP PPPTPTP   PPT P T                      T        TP   PTPPPPP  PPPP  PTPPPTPPPP T   TT T T                      T   T          T           T   T      T                   PP  PPP   PT PPP    PPPTPPPPPPPPT  TTP  PPPPPPT  PP  PPTPTTTPT    PP PPP PPP PPPPPPPPPPPP T TPPPPPPP TPPPPP PP  PPPP PP  P  PPP PP TPTTPP  P TPPP PPPPPP PTPPPPP T    P   PPP PPPTTPP TTTPPPPPTP   TTPPTPTPPP  TP   P PPPPT T PTPPPPPTPP PPPPP PT TT      T    T T           TT   PPP P PPP  P   PPPPPT  PPPP PPPTPPPTP P P   PPP TPPP PPT TPPPTPP PT  TPPP PTPP    PP PP PP  PPPPP PPTPPPPTPPPP TPP  TPP PPPP   PPP PPP TPPTPT  P PPPTPPP                     T      T   TPPT PPP PPTPTP P PPT P PP PPTTPPPP  PP PPPPPPPPP  PTPPP  T P   PPTPPPPP  PPPPPTP P PTP   PPP PPPP T T    PPPP PP PP  P TPP PPP PPPPPPTPPPPPPPPPPPP PPPPPPP P PPPPPPP TPP P TT  P TPTTPPP PPPP PPTPPPP PP PPTPTPPTPPP  PTPPPP T   PPPTPPP PPPPP P PPPP  PP P PP  PP PPPTPPPPPPP   T PPPPPPPPPPT TPPPP PPPPPPP  PP  PPP  PTP   P  PPTP  PPP PPP  PPPTTPPTT  PPT  TPP TPPPP TPPP PPPPPPPT     P PP  TPPP  P TPPP  TTTPPPPP   PPPPPPT P TPP PPPP  PP  PPPPPP PPPPPT TPPPPPP TP  PPPPPPTP    PP PTPPPTTPTPPPPTPPPPPPP   PP  PPP  PP P PPPPPPPP P PTTPPPTTTTPTPT P P PT    T                         PPPPTPPPPPPPP P  PPPP PPPT PPPP TPPT TPPP  TPPTPPPPPPPTPPPPPPPPPPPPPPPPPP  TPTPPPPPTPPPT                        T         PPPP  PPPPTTTTPTTT PP  P  T TP             T            T  TPPPPPPT   PPP PP   TTPPPPPPP  PTPPP TPPPPPT  P  P  PTTP  PP  P     PP PPPPPP PPPPPP  PPTP          T     T      TT       PPTPP P  PPPP  PPPPPT PP PPPT P P   P  TPPPPP   PPP PPPPP PPPPT PPPP   T  PPPTT    PPT   PPP PTPPPPPPPPPPPTTPTPPPTP  TPPPPPPPPTT PPPPP  PPPPPPPP PPP TPPPPPPPPPPPPP PTPPT TTPPPP  T  PPP PPPP P T  PPPPPPP  P PPPPPP  TPP     P  PPPPPPPPPTTPP P  PP    PP PTP PPPP PPPP PPPPPTPPPP T  PPPPPPTPP PPP  PPPT  PP  TPPPTPP    PPPPPPPPPPPPP PPPP TPPT PP P   TPPT PP PPPPPP PPPPPPPT PPPPP        PPPTPPPT P PPP P P PPPPPPPTPPP    TPPP TPPPP  PP TTPTPPPPPP  PPPPPPPPPP P PPP  PPPPPPPPP PPPPPPP PP  PPPTPP  PPPPPPTPP    TPPTTPT PPPP PPPP  P  PTPPPPPP PPPPPP PPPPPPPTPPPTP     PP  PPP PTP      PPPTTPTP PPTPTPPPPTP  PP    PPP  P TPT TP PPT PT P PP P TPP        T            T TT       P  P  PPTP PPPP T  PPPPTTPPPPPP PT T T  T TP PPPP PPT PT     PPTP P PPPP PPT  PPPPPPT  TPPTP PTPPPTP  PPT  PPPPPPP   TPPPPT  PPPP   PT PP   T    PPP  PTT T      T          T         P PP PPPPPPP PPP PTPPP  TPPPPPPPPPTP PTTTPTT PPP PPP TPP  PPPPPP P TP P PTP   TP  PPPP PPPTP TTT    TPPP PTPTPPPP  PP  P PP  PPT PTPPP TPTPPP  PT P  PP        T    T   T   T    T     PP TT PPP  TTP   T PPTP P PPPP   PPPPPT TPT  PP PPT P TTP TPPPPPPTTPTP  PPPPP  PPPTPPPTPPP PPPTPPT PPT TP PPPPPTPP  P   T        T T             T   T PPP P   TPPP  T  PPPT TPPP P                   T TT          PP P TTP  TTPPPPPPPTTP PT     PP PPPTTTTPPPP PP  PTPPT PP PP PPPPP    PPT TP PP     PTPPTPPPPPTT PPT PPP  P PPPTT PP  PPPPP T  PT    PPTPT  P   TP  P  TTT  T   T TT TTPPP T     T  PTT    PP TP TTP PPP P PPPPPP   PTTP PT   PPPTTTT  T PPPPP P TPPPTPT   PP PP T PPT T   PPPPTPPP  P TPP PP  TPP     PPPT P P T      T            T      T                       T     T    PTTT  PPP   T   P PP  PTP  PT  T  T  T  T   TTTT   T      P  P   P PT TP     TPPTPPP PPP PPT PP P PPP   T  PPPPPPPP PPTP P PPPT    PPP   T  P PP  PPTP  PT  P   T TT PPPPT PPP PTPPPT  PPPTPPPPP PPPP PPPPPPP PPPPPPP PPPPP P   TPP  PPPT  PT P  P   PPPPP  TPPPPPP PPP P     PPPPP   PPPPPPPP  PPPT PPP TP  PPP PPPPP  PP PPPP    PP  PPP   PPPPPT   PPPPPT  PPPPP P PPPTPTTPT PT  PPT PTTPPPPPPP  TPPPPP  PP  PP    PP  P  PPPPPPP PT    PPP     PPT P         PPP    PPP PT   PPP T  PP      PPPPPPP PP TPTP    PTPT PPP TPPPPPPTPP   P TTPTT TPPTP  PPT   PPPPPPP P P PPT  P   PP   PP   PPPPT PP  PP PPT  T  TTTPPPPT P  T P TPPPPP P  PT P TPPPP TPPP  PPPPP   P    PPP PPP      P  TPPPP  TPPPPT PPP PTPPPPPPPT PP  T T               TT        PPTPPTPPTPP   TP PT TPPPPP   PPPPPT  TTPPPPPT   PPTT   PP PPT            T T   T            PPTPPP PTTT  PPPPP  P   TPTTPP    PPP PTT P   P PPPTP PPTP P  PPPP   PPPPPPP  PT PPPPPPT  PPT PPT P  P   P  TP  T    TPPPP  TTPTPPP   PPP  TP    P   PT  PPPPPTPP P TPP          PP        T  TT      T             PTTPPT PPT TT T     PTPPPPT  PPPPPT PPPPPP  PPPPP P   PP  TPPPPT  P  PPPPPPP T  PT   P PPP  T        T     T   TT    T  PPPPT PPP PP  PTP  P  P TTTPT  P   PP PP  PPP  PPP P PPP P  PP   PPTP   P  PPT P PPP P P PT PPP  P  P PP     PP PPP     TP PPPPPTTTT  PPPPPPT  PPPPTTPPT PTPPPP T P  PPP   PP PPPPT   PPPTTTP TPPT PPP PTP P PPT  TTPPPPPPP PPPPP  TPT TPPP    T   P TP P  P PP PPPPPP PPPPPP TPT   TP PPPPPTPPPPPPPP  PPTT  P   PPP  PPPPPPPPPPPP    PPPTPPPTT  PP PTPPTP  PPPPP TPPPPP T  TPPPPTTP PPT    PTT PPPP PPPPPPPP T P   P  PP  PP    PPTTP  PP   TT PPPPPP   PP P   PPPPPPP TP   PP  PP   P      TPPTT PPPTP TPPTP PTPPPP  PPP   TPP  P    PPPPPTT TPTPTPPTTPPPTTT PT P P   PPP PP  PPT  PPPP TPPPT PPTPPPPT TPPPT T     PPPP         PPPPPPP   PP PPPPPPP PP  PPPPT TPPPP  PPPPPTTPPT PPPT PP T PP  PP PTPP     TTPPPPPP P  TTP PTP PP PPPP  P  PPPPPPPP T   PP   PPPPTPPPPP     PPP   T  PPTPPTPPP  PPPPP    PPPTTTPPPP  PTTPP   P P PPTTPPPPPP  PPPPTP  PP  PPPPPPPPPPPTPPPPP PPPPPPPTPPPTP   PPPPT   PPPP  PPPP  T  P   PPPPPT P TTPPPPPTTPPPPPTPP      PP  T PP TP PPPPPPPT  PPPPPPPPPPPP PPP PP  PPPP PTPPPPPPPTTTPPPPTPPPPPPPPPPPPPPPPPPPP  PPPPPP PPPPT PT PPPTP PP PP   PPT  PPPPPPPPPPPPPTP  PPPPPPPTPT  PPPPPP  PPPPP PP  PTPPPPP  P PPPTP P PPPPPP  TPPPP P  P  PP  T TPPPPPPP  PTPPPPPPPPT T  P PP PTPP PT  TP  TPPPPT   PPPPPPPP   PPPPPTTPTPPPPPPPP PPPPTPP  TPPPPPT  PPPP TPPPTPPPPT PTT P PPT  TPP PTPTT PPT  PP  PPPPTPPP PPPPPT PT PPT   T    PTT T    T   PT  PPPP  PPPP PPPPPPPP TTTP  PPP  P PPPPP   PPPPPP  PPPPPP      PP T     PPPP P PPTTTT  PPPPPPTPP     PTPT T PPP PP PPP PP P P PP PP P    T T PPP PP PPPPPT  PPPPPTT       P    PPT   TPPPPPPTPPT   PPP PP  PPPT  PP  P  T TPPPP PPPP TP PP P P P PP P   TPPPPPPP  P PPPPT  T T P PPPT  PP  PT     PPPPPP PPPP PPP PP PP PPP   PPPPTPPPPP PP P  PPPPPPPPPP P PPP TPP TP PPPPPP PP   P PPPPP   PPPPPPPPPPPP   PPPP PP     TPPP PP P  P PTPPPPPPPP PPPPPPPPPPP PP P  TPPPPPPPPPPPPPP  PPPPPP    PPTPPPPP  PPPPTP PPPP PPP P PPPPP P  PT P  PPP  PP  P  PP  P  PPP  PPP    TP  PP P   P  T  P PPT PP  PP P T   P  PPPPPPPP PPPPPPTPPTPP  PT  PP PPPPTPPPP PP  PP  PPPT  PP  PPPP PPPPPPPPPPPPT PP PP  PPPP P P P   PPT  PPPPPPPPPTPPP P PPPT PPP PPPP PPPP    PP   P PPPPPP   P  PPP P PP  PPPPP   PPPP  PPP               T       T      PTPPPPP TP  TPPPPP PP PP T  P   TPPPP   P       PPTP  TPTPP PPPPPP PP PPPP  P   PP   PP P  T  T   PP P P  PPPP   PPPPPP     T PPPPP TP     PT PP    PPP    PPP P  PP PP   PPP PP    PPPP PTPPPP  PPPPPP   P PPP PP PP  P   PPTPPP       P   PP    T PP P TPPPPPPPTPPPPPPP    PPPPPP PPPPPPTP PPP     PPP TPPT P   PPP  P PPPPPPPPPPPP      PPPPPPP PPP TP     PPT  P TTPPP   PP     PP TPP TPPP PP PP  P    PPPPPT P  P PPPPPPPT PPT P PP  PPTPT  P T PT TPPP  PPPT PT PTTPPPP  PPPPP PP  PPPP    P  PPT TPPP  PP PPPTPPPPPPPT   P P  P  PP PPT    PP  T PPPPT   PPP   PTPPPPPTT  PP    TPPPPPP      T  PPPP  P PPPPPP   P PPPPPTPTPP  PPPPP PP    PPP PP PPP  PP PPP  PPPPPPPPPPPP PT  PP   PPPPPPPP     PPPP P  PPPP T PPPPP TPPP PP  PPPP  PPP PPPTTPPPPPPPPPPPPPP  PTPP P  PPPPPP        T  PPPP P    PP PPPPP  PPP PPPP PP PPPPPPPPPPP  PPPPPPPP    TP  PP P   TPPP  PPP PTPP T      PPPPP PP      T   PPP PPPTPPP   PPPP   P PPPPPP      P  P P   P P P PPP     PPPP PPP PPPPPP  PPPPPPP PP  PPPP    PPPP      PPPPPP P PPPP P  PPPPPPPPPPP  PPPPPPP   PPPPPPPPP  T  P  P P PP  PP  PPPPP    PPPPPPPPP PP T  PPPP PPPPPP PP PPPPP   P   P PP  PPP   P     PTPPPPPPP   T PP    PP PPPP P P P PP   PP P   PPPP  P  PP  PP  PPP  TPPTP PPT  P PPPPPPPP  PP TP                                T  T    T  TT                       T         T          T       T   T                        T    T   T                                    T     T  T  T      TT  T  TT              TT          T           T       T       T      T T   T     T                    T    TT            T                                             T T   T                      ", "T    T  T         T T T    T      TT            T  TT                T                            T         T          T   T T   T                     T           T           TT           T    T           TT   TTT      T      T           T      T   T                   T T                       TT               T             T      T    T    T T               T    T  T T  T  T      TT                T        T TT     T                T  T                            T      T T T                                               T     TT                 TT  TT   T              T    T      T                               T   T                     TT  T  T   T     T        T  T              T            T                       T              T           T   T       T              T                                        T T              T T  T        T              T T    T      T     TT                                       T        T       T            T       T                        T                        T        T            T  T     TTT   T         T            T T    T       T                             T                                         T          T                                      T           T                          T                                        TT T T                    TT           T           T                                  TT                     T      T T T           TT          TT                        T          T    T        T             T                                   T                          T                   T                          T                 T            T  TT       T         T            T T     T       T      T TT  T     TT     T    T               T T                         T       T               T   T             T   T       T                         T    T        T    T                                                   TT                   T        T                                     T           T T                     T T   TT   T                                  T    T   T                               T     T         T   T T        T          T                   T              T         TT  T   T   T        T T     T                                                      T   T                        T  T                    T TT T         T            T           T       T             T          T               T           T    T        T   TTT     T  T          TT    T               T T  T                                                                                                                     TT                                                            TT                    T                                                                 TT  T               T      T  TT         T T                      TT                                                                                                         T        T                             T                                                  T                                                                                 T                                          T               T        T      T                                   T                                                      T                        T    T                    T  T                 T             T                T      T              T   T                 T   T      T                       TT                        T              T      T           T                   T    T  T                                       T                         T                       T T                        T                                   T               T             T                                            T      T                                      T   T   T       T         T   T                                                   T       T  T T                                                                                  T         T T                                                                                                                        T            T                                T          T    T                                                     T         T                 T                                  T                   T              T                                                                    T    T                                          T                                        T                           T                                                              T         T       TT   T                                           T        T   T                          T                                                                      T     T                   T       T                        T            T              T              T     T     T                            T                                 T           T                         T TT                              T                                                                     T    T      T                                                                                        T                   T               T        T     T                                       T      TT             T T                           T  T TT T        T      T     T                 T  T            T  T  T  TT          T            T              T      T               T                       T            T T                  T                                                       T   T                                        T                 T  T T                    T               T                    T                       T     T               T T   T       T          TT                     T T                                          T    T            T                       T                       T                                        T                                                T                       T        TT    T               T  T    T                      T     T TT               T                T                     T    T             T T                                                                                                       TT                                         T                                            T                  T      TT         T                            T      T       T          T T   TT     T                                                                                                                  TT  T                                    T                                                                                     T  T         T   T         T                  T      T           T    TT                                      T                     T   T                                                         T                                 T                        T                               T                                                                T              T      T T T   T  T       T  T       T                         T        T                     T   TT         T     T                   T     T          T  T                                               T                            T             T       T             T                                  T            T                                         T            T       T            T     TT       T T  T T        T  T TT TT        T                     T                           T             T   T           T                                        T         T           T     T       T             T   T            T     T T                                                                                                         T       T               T            T                    T       T                      T     T        T                                                                                          T                      T                T  T                         ", "                                      T                     T         T                                           TT                             T                            T                        T TT T                 T                                             TT                                     T T                     T      TT                   T                         T                             T         T T        T T                      T                                  T                                   T       T         T  T         T  TT    T  T                                       T       T                             T                                                                     T T T                                                           T       T             T        T                             T             T   T   T T T     T                               T                     T   T                                     T                                                                                  T           T           T                                            T                             T                                      T                                                         T       T                    T                       T                              T                                                                         T                                       T     T         T   T   T                             T              T           T       T       TT                            T       T              T                 T T                          T                     T                        TT            T                                                                                                                                                            T          T                              TT          T       TT     T T              T              T T   TT   T                                                          T        TT   T                 T      T                 T                             T             T     T                                   T        T T            T   T       T                                                        T                                                                                                           T                                                              T           T                            T                                                                                                                T T                       T      TT                     T                                                                                        T T    T                      T            T                                                                                    TT                                       T                                 T                        TT                     T               T              TT              T                                                 T                       T                                                                                                                           T      TT            T             T                       T   T                                T            T  T                   T                            T                 T             T              T                  T                                           T                                                           TTT                              T       T    T                  T                        T          T T T     TTT              T     T   T                    T                               T      T                                                          T          T   T         TT                                                                            T                                                                 T                   T                             T       P                          P              T               P             T                                                                                                           P                              T                                   T      T                      T             T                                 T                                       PPP                                                                                         T                   T                                                                      T                                                     T                                                                                T   T     T                       TT                T                     T                                                                                                                                                                                                                                                         T               P                                                     TT               TT T     T     T      T  T T                                                                        P                                                                                                                                                                                      T                                                                          T                                                                                                                                        T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    T T     T                                                                        T              T                                                                                                                                                                                                                                           T                                       T                   T                                                                                                                                                                                           T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                T                                                                         T T             T                 T                                                         T                             T                   T       T         T                                                                                                          T   T                                                                                      T           T           T T                     T                           P                    T              T            TT                                                                             T                           T        T                     T  T      T                  T         T   T                                                      ", "         T                                      T                                   T                  T                                        T                                           T                                                  T   T T                    T                     T                                       T                                              T  T                        T                                                                                          T     T                     T       T      T                                     T                      T              T    T                   T                T                                        T          T                   T                        T  T                                     T       T                     T             T                                                 T    T        T                                                                                TT                                             T                 T                                                                         T   T            T              T T                                    T T  T                                               T  T                                       T                        T                                               T       T   T           T                   T                     T                                                                       T                            T                                     T            T                                                                                   T                                            T           T                                                                                T       TT         T                        T         T                        T               T                                      TT                                                                                  T                                          T                                                                                                  T     T           T                                                                            T                                                                        T        T    T                                     T                                                T                                          PPPPPPPPP   P P   P P PPPPPPP PPPPP PP  PPPPP  P    PPPPPPPP P                           T                 T   T      T TT    TT             T                            T             T            T    T                                                                                                                                                            T                   T                                                        T                TP           T      T  T       T      T       T                        T                                                                                                                                                    T               T                                T                                           T        T                                 T                                                                           T    T        T         T          T                                                  T         T      T  T         T                T                   T                 T  T                                                                    T                                                                 T                T            T                                         T                                                           T    T    T                          T                                T                                    T                  T             T      T                        T            T    T                     T                                                                T                            T                            T          T                                                                                                                                         T            T   T                                                                    T                    T    T      T                       T                                     T        T                    T                                                 T                                                                         T                                                                            TT                                                                                                        T                                                T                                                                                                                                                             T                                  T         T                               T      T    T                                                                    T         T                              T   T       T                                              T  T                                                             T        T                       T                      T        T                T            P  PP  TPP PP   PPP    PPPPP T T      PTTPPP   PPPPPPP        P          P PTT    T TPPPTPP  PPPPPPPPPPP PPTPPPP  P   TP P  PPP TPT P  TPPPP TPP PPPP  TTPPPPPPPT     PP  TPPPP   P P TPP PPT PPPPPPP    PTPPP PP  P   PTPPPPPPP    PPPP  PP   PTPP    P  P  PPP   PP   PPPP  PPPP                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              T        T                  T   T T                                      T       T       T      T T                                                       T              T               T  T     T                               T                                      T           T       T         T          T            T                          T                                    T       T T                             T          TT                             T      T                       T  T  T  T       T      TT          T  T                T                   T                            T                                                    T                                 T                                                           T                                T                                           T  T                                  T                 T   T        TT       T  T                                                 T                     T       T                   T          T         T                  T      T                                            T T                T                                 T                  T  T                                                            T                                                                                     T                                    T T     T    T                                                  T T    T                T     T  TT             T    T               T           T      T                                                                      T           T   T                             T                                 T ", "                                                                                T    T   T                         T                                       T                                 T      T                  T                     T            TT       T                 T                    T                                                                                                                                                                             T         T                       T       T                   T     T   T                                                      TT    T                                                        T                                                    T                                                                         T                                        T             T                                                            TTT                                        PP                        T                                                                                                  T          T     T         T             T                                           T                                                    T                                                          T                               T            T  T         T               T            T                                         T                 T          T T    T          T                                                                  T          T                                                  T       T                     T                         TT           T       T                                                             T       T         T                                   T        T                                   T        T                       T T                                                                         T                        T                                              T                                                     T                          T       T                                T                     PP                                                        T             T                        T T                   T                      T               TT  T   T     T                                                                              T                                        T                                     T                      T    T    TTT     T                                                   T                                      T    T                                                                                                                    T  T                                                   T                                                   T              T            T                T                                                 T                T            T                 T        T                      T                      T                                    T           T             T              T T      T                                                                          T                            T                                 T           T                     T        T                                                                     T                                               T              T     T                T      T           T      T                                       T        TT T   T                                                  T     T   T                                         T                        T                                  T   T                                                  PPPPPPPPPP  P     P   TPPPPP  P       T                                    TT            T         T                                       T T                     T   T      T                             T                                                                                                                               T              T                         P                     TT   T               T      T                     T   T                  T    T     T              T                                                             T                                               T                         T  T                              T        T                                               T              T       T      T                T T               T               T                             T    T   T    T                                                 T                                                                         T  T                                      T       T                                                                                        T        TT                          T                                     T                                                           T        T                                                                  T    T                                                         T              T                                                                 T  T          T     T                        T                              T                                  T                                        T                                                            T  T                                                                                  P               T P                     T                T   T                              TP                                                T                                                           T                 T   T        T                           T                  T                    T  T                                     T                         P        T                              T                                           T                 T                P               T                   TT           T                    T      TT              T T      T                      TT    T                    P                                       T                        TT                                  T                T      T  P   TT          T             T   T         T              T T                   T T                               TP       T                                          T    TT                          T                                                                                                                                    T                 T                                           T                     T        T                      T                             T      T                                                                     T      T        T                T   TT                  T                                                                    T      T   T   T  T                                                                           T                           T                                                         T                                    T    TT                             T PPP  PPPPPPP PP  PPP P PPP   PP   T                          P  PPP P PPT PPPP PPPPPPP PPPPPPPP P PPPPPPP PPPPPPPP PPPP PPPPPPPPPPP PPPPP PPPPP PPPPP PPP                 T            PPPPPP PPP PPP PTP P PP P  PP PPPP PPPP PPP P PPPPPP PP  PP                               PP PPP PPP PPPPPPPP  PPPP P P                                                                                           PPPPP PP  PPPPPP    PPPPPP   P                                                                                           P PPPPP P P PPP PPPP PPPP PP PPP PPPPP PPPPPPPTPPPPTPTPPPP P PPPPP  PP PPP PPPPPPP  PPPPPP   PPPPP PPP PPPPPPPPPPPPPP P  P  P PPPPPPP PPP PPP PPP  PPPPPPPP PPP TTPPPTPPPPPP P PP PP  PPP  PPPP PPP PPPPPPPPP P PPPPPPP P  PPP PPP   PP PPPPPPPP P PPPPP PPPPPPPPPPT  PPPPPPPPPPPPPPPPPP PPP  PPPPPPPPPPPPPPPPP PPPPPPPPPPPPPP PPPPPPPPPP PPPPPPPPPPP PPP PPPPPPPPPPPPP P P ", "P                T T   T        PPPPPPPPP TPPP PP PPPP P  PP P PPPPPPPP PPPPPPPP PPPP PPPPPPP  PPPPPPPPPP PPP    PPPPPP PP PPPPPPP P PPP P  P P PPP PP PPPP PP     PPPP P PPP  P PP P PPPPPPPPPPPPPP  PPP PP PP PPPPPP PPPPP PPPP P PPPPPPPPPPPPPPPP PPP PPPPPPP PPPPPPPPPPP PPPPPPPTPPP PPPPP P PPPPPPPP PPPPPPP PPPPPPPP PPPPPP PPPPPPPPPPPPP P                                                                                        PPPPP PP PPPPP P PPPPPPPP PPPPP  P PPPPPP P PPPPPPPPPPPPPP   PPPP PP PPPP PP  PP PPP PPPPPPPPPPPP PPP P PPPP  PP PPPPP  PP                                                             P PPPPPPPPPPPPPPPPP PP PP  P PP                               PPPPP PPP P PPP PP PPP PPPPPPP PPPPPPPPPPPPPPPPPPP PPPPPTPP                              PPPP PPPPP PPP PPPPPPPP P P PPPPPPPP PPP P P  PPPPPP  P PPPPPPPPPPPPPPP PPPPPPP P  PPPPP PPPPPPP PPPPPP PPPPP P PPPP   PPPPPPPPPP  P  PPPPP PPPPPPPPPPPPPPPPPPP PPPPPPPP PTPPPP PPPPPPPPPPP PPPPP PP PPPP PP PPP PPP PPPPP PPP PP PPPPP PPP PP PPP PPPP PPPPPPPPPPPP PP P PPPPPPPPP                               PP P   PPPPP PP P PPPPPPPP P                              PPPPPP  PP P PPP  PPPPPPPPPPPPP                              PPPPP P PPPP P   PPPPPP P PPPPPP PPP PPPP PP  PPP P PPPPPPPP P                                                              P PPPP PP PPPPPPPPPP PPPPPPPP                              PPPPPPPPPPP PPPPP P PPPPP P PPPPPPP PP PP P PPPPPP PPPP PPP PPPPTPPPP PPP PPP TPPPPP PPPP PPPPPPPPPPPP PPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPP PPPPP PPPPPPTPPPPPP PPPPP  P PPPPPPPPPPPPP                 T            PPPPPP PPPPPPP  PPPPPPPPPPPPPPP   T                                                         P PPPP PPPPPPPPPPPPPPPP PPPPP                           T                                PP PPPPPPPPPPPPPPPPPPP PPPPP                              PP PPP PPPPPP  PPPPPPPPPPPPPPP                                                            PP PPPPPPP PPPPPP PPPPPPPPPP P                              PPPP PPPPP PPPPPPPPPPPP PPPP P                  T           PPPPPPPPPPPPPPPPP PPP PPPP PPP P PPPPPPPPPPPPPP PPPP PPP PPP PP PPP PPPTPPPPPPPPPPPPPP P T                              PP PPPP PPPP PPPPPP PPPP P PPPP                              PP P  PPPPPPPPPPP P  PP  PPPPPP               T     T        P P PPPP PPTTPPPPPP P P     P PPPP PPPPP  PPPPPPPPPPPPPP  PPPPPPP PPPTPPP PP PPPP PPP PPP PPP P P TPPP PPPPPPPP PPP PP PP P                            PPPPPPTP P PPPPPPPPPPP PPPPPP P                                    T                  T    PPPPP  PP    T PPPPT P  PPTP P   T                                                         PPPPP P P PPPPP   PPPPPPPPPPPP                              PPPP  PPPPPPP P   PPPPPTPPPP PP  PPPPP   P PPPPPP PPP   PPPTPP  PPPP PP   PP PPPTP  PP PP  PTPPPPPTPPPPPPP PPP PP PPPP   PP PPP  PP  P  PP PP  PPP  PPP  PPPPPPP  P PPPPPPTPPPPPP   PPPPPPPPPPP PPPP PP PPPPPPPPPPPP        T                        PPP   P PP PP  PPPP P  P  PPPP PPP PPP PPPPP PP PPP PPPPPPPPP PPPPPPPPPPPP PPPPTPPPPPP PPPPPPPPTPPPPP PPPPPPPP PPPP PPPPPPPPPP PP   P  PPPPPPPP PPP PP PP P  PPP   PP  P PPPPP    PPPPP   P  PPPP P PPPPPPPPP   PPP P PPPT PT PP  PPPPPP PP PT PTTPPPPP    PPPPPPPPP   PT P PP PPPPP  PPPPP     PPPPP PP T TP PPPP P PPPPPPP  P PPPP PPP PPP  PPP P  PPP PPPPPP PP   PTPPPPP  P P PPP    PPPPP P    PTP  PTP TP P   P PT PPPPPP PP  PPPPP            T                 PP PPPPPPPT PPPPPPP PPPP  PPPPPPPPPP PPPPPPPPPTPP  PPPPTPPP  PP PPPPP  PPPP   PPP P PPPPP PP P  PPPP PPP    P PPPPP PP  PPPPPPP PP  PPP P PPTPP  PP P          TT                  T   PPPP PP   PPP PPPPP   PPPPPPTPPPPPP P PPPPPPPPPPPPPPPPP   PP  PPP PPP  P PPP   PP   P   PPPP  PPPP T  PP    PPP   PPPP  P   PPPPP P    PPP PPP PP     PPPP PPPPPPP  P  PPPPPPP PPP P   PP   PP  PPPPP PP     P PPPPP  PPPPPPPPP PPP  PP  PPPPPPPPPPPPPPP PPTP PPPPP      PPPPP P   PP PPP  PP P      PPPPP  P P P  P  PPTPPPPPPPPPP   PP  P PP PPT P P  P P PP   P PPPPPPPP                                 P P    P PPPP  P  PPT    PPP   PP  P PP  T PPPP PPPPPP PP  P PPPP TPPP PPPPTT PPPPP PPP PPPPP P PP  PPTPPP  P P P PPPPPPPPP  P P T   PPPPPPTPP  PPPP  P PP  PP PPPTPPPPPPP  PPPPPP  PPP  PP  P  PP PPPP  P      PPPP  P  PPP  PPP  PPPPPPP PPPPPP  PPP  P  PPP   P PPPPPP  PP P PP PPPT PPPPPP   PTP  PP PP PPP  PPP PP PPPPPP P  TPP PPPPP T T PPP P P  PPP  P  PPPPPPP TP   P      TPPPP PPP P   PPPPPP   PP PPPPPP PPPP PPPPPPPPTPPPPP P PPPPPPP P   PPPPPP      PPP  PPP  T  PP PPTPPP PPTPP    PPPP PPP PPPP PPPPPPPPPPPPPPPP  PPPPPPPPPP  PPPPPPPPPPP        PPPPTPPPPPPP P  PP PPPPPPPP PPPPPP  P PPP  PPPP  PPP  P  PPPP             T                TTPPPPP T P PP PP  P  P    PP P   P  P PPP  PPTP PPPP   P P  P  PPPPP TPPP  PPPP    PPP   P PPPPPP P  PPPPPPPPP   PP   PPTPP    P    P   PP PPPPPPP   PPP PPP  PPPPPP P  P PP   PPTPPPP PT PP PPPPPPPP  PPPPPPPPPPP PPPPP  PPPP PPPPPP PPPP     P PPPPPPPPPPPPP PT PP  P  P PPPPPPPP   P PP PPPPPPP PPPPP    PPPPPPTPPP  PPPT  PTPPPPPPPP  TP PPPPPPT  PPPPPP  PP  P  PP  TT PP P PP PP  P PPPPP PP  PPPPP    PPP PP     TPPPPPPPPPPPPPPPPPPP P PPTPPTPPPP   P  P   PPP PP PPPP  P  PTPPP PP P P  PPPT                               PPP PP  PP   TPT  PPPPPPPPPPPT P PP PP    PP      PPTPTPP P PP   TPP PPPPPPPPPPPPTPPPPPPPTPPPPPPPP   PPPPPPPPP    PP PP PPPPP   PPPPPPPPP PPPPPP PP  P  PPPPT   PPP TPPPPP  PPPP  PPPT P        T                       T      T   T              PTPTP T P PP    PP  PPTPPP    PPP   PT   PPP  PPP  P  PPPPPPTP PPPPP PTPP PPPTPPPPPTPPPPPPPP PPT  P PPPP   TT PPPPP P P PPPPPPPP  P TPP PP PP   P   PPPPPPP   PPPP P P   P PPPPPT    T   PP PPPPPP TPP PPPPP  PPPPPP  P  PPP PPP PPP PP  P P PPPPPPPPPPPP   P  PP P PP PP PP  PP  PPPP PPPPPPPPPT   PPPP      PPP  PTPPP   PP TP PPP PPPP P  P  TT P PPPPPPPPTP  PP    PP   PP PP T  TPPP  P PPP P  P  PPP  PP  PPPT PPPP  P   PPP  PPP P  PPPPP   PPP PP   PPPPPTPPPPP PP                              PPPPPPPPPPP PP PP  P  P   PP TP   PPPPPTTPPP PPP    TPPPPPP PP PP PP PPPP PTP P   PPP    PPP                  T             PPP  PPPPP PPPPPPPP PPPPP PPPP    PTPP PPPPPP  PPPP PP PP PPP PPP  TP  PPP T PP P   P PPPP P  PPPPPP PPPPP PPP  PTTP  P PPPTPPPT P    PPP  PPPP  PPP PP P TPPPPP      PPPPP  PP   P                              PPP PP  PPPPPPPPPPPP    PPP PPPP PP PP PPP PPPP PP PP PPPPPPPT PPPP PPP   TPPP  PPP PPP P PPP PPPP  PPPPPPPP      PPPPPPPP            T                 PPPPPPP PPPPP   PPPPPPPPP   PP   PPP  PPTPPPPPPPPPPP    PPPPPPP  PPPPPPPTPPPPPPPP PP  PPPPP PPPTP  PPP P  P PP   P  PPPP  PP   PPP PPPPPP P P PPP P P P P PPPPP PPPPP  PPP PPPP  PPP PPPP PP  PPPP PPPPPPPPTPPPP PPP        T    T                PTPPPT PPPP  PPP    PP   PPPPP                           T PPPPP  PPPPPPPPPPPT PPPPPPPPPPPPP  P PPPP   PPPPPPPTPPPPP TPPPPP PPPPPPP  PP  PP  P    PP  PP   PTPPPPPP  P  PP    PPPPPP   P  PP  PP PPP  PP   PPPPPP PP     P  P P  P  TPPPTPPPPPP   PP PPPP TPPPPPPPPPT P PPPPPPPPP                              PPPPTPPPPPPTP  PPP PPPPTPPPPPPP PPPPPT PPP PPP  PPPPPPP PP PPT PPP  PP P  PP TPPPPP PPPPPP P   PPPPP  PP  PP PPPPPP TPTPTP   P P PT PPP PPPPP   PPPP PPPPP  PPP  PP P PP PPPP  P P PPPPPPP   P PPPP P  PPPPP  P PP   PP  PP PP  PPPP   TP  PP PPPPPPPPPPPPPT PPPTTPPPT   P   PTPPPPPPPPPPPTPPP PP PPPP PPPPPP PPPPPPPP  P PPPPP PPP PPPTTPPPP  PPPPPPPPPPPP  PT P  PPPPPPPPPPP PPPTPPPP P    PPPPPPP  PPPP  PPPP PPP P  P  PPP PP PPPP  PPPTP P  PPPPPPP P PPPP  PP PP  TP PPP PPP PPPPP  PPP P   PPT      PP PP PP  P PPP  P PP  TPPPPPP   P PPP PPPPPPPP PPP  PPP  P   P  PPTPPPPPPP PP PPP   PPPPPPP  P    P  PPPPPPPPPPPPP  PP PPPP    P   P       PPPPPPPPPPTPPPPP PPPPP  PPPP P   PPPT   PPPP P PPPPPP  PPPPPPPPPPP PPPPPPP PP P   PPPP P PPP PP  P PPPPPPPPPPPPPPPPPPPPPP PPPTP P  PPPPPP  TP    P PPPPPPP  PP PP       T                       PPPPTP P PPPPP PPP  P  PP PPTPPP P PTPP    PPPPP  PP PPPPPPPP PPPPP     PPPP  P PPP PPPP  PP  PPPPP PP PPPPPPP PTPPPPPP PP PPP PPPP P PPPPPPP PPP PPP  PPPP PPPPTPPPPP P PPPPPPP PP   PPPTPPPP PP P PPPPPPPPPPPPP TP PPPPT  PPPPPPPPP P  PPPP  PPP PPPP PPPPP P PPPPP PPPPPPPPPP PPPPPPPPPPPPPPPP   PPPPPPPP  PP  PTPPPP   P   PPPPP   P PPPPP   PP PPPPPPPP P  PPPP  P PPPPP         T  T                PPP  PP P PP P P    PPP", "PP  PPP PPP PPPPP  TP    PPPPP PPPPPP  PPP      PPP P PPPPTP  PPPPPPPPPPP P  PPPPPPPPPPPPPPPP   PPPPPPPP PP  P P         PPPPPTPPPPPP    PPPP   P P  PPPP PP P   PPPPPPPPPP PPPPPPPPPP  PPPPPP PPPPTPPP P     PPPPPP    PPPPPP    PPPPP   PPPPPPPP P P TPT PPPPP     P T PP P TPPP PPPP TP PTPPPT  PPPPPP  P PP    P PPPPTPP   PPP PP P PPPPPP PT PPP PPPT  TPPPP   P  P  PPPPP  P PP       T           TT          PPPPP  PPPT   PPPPP  PTP PPPPPPP   PPPPPT T P   PP PT PPPPPPPP PPPP PPP  P PP  PPPPP PPPPPP  PP   PPP   TP      P  T P PPPPPPPP PP  PPPPPPPPPPPPPPPPPTP  PPPPPPPPPPPPPPPPPTPPPPPPPP PPPPP PPPPP P  PP   PPPP  PPP  PP PPP PPPPTPPP PTTPPPP  PPP  PPPPPPPPPP P   P  PPPPPPPPPPPPPPP   PPP PP T PPPPPPPP    PPP                                                                     PPPPT   P PPPPPPPP  PP  PPPPPPPT PPP PPPP  PPPPT PTTPP   PPPPPP T P    PPP PPPP PPP   P   PPP PPPP   P PPPPPPPPPPPTPPPPPPPP PPTP PPPPPPPP  PPPP PP PP PPPP PPP PPPPPPP PPPPPPPPPP   PPPPPP  P P PPTPP  PP P P  PP    PPPTPPT  PPP PPPP P PPPTPPPPP  PPP P PPPPT     PPPPPP  PPP PP T PT    P  PP P PPPPP PP P PP  P  PPP PPPP  PPPPPP P   PPTPP PPP  P  PP    PPPPPPPPPPP    PPPPP PP P   PPTPPPT PPPP                              P    PP PPPPP PPP   PPPPPP P PP  PTP   PPP   PPPP PPPPP P  PP   P PPPTPPT PPPPPPPPPPPPPPPPPPPPPPPP    PPPP   PPPPPP PPPPPPPPPTPPP PPPPPPP  PPTPPPPPPPTPPPPT P P  P P P  P PPPPPPPPPP  PP P  PPP  PPPPP PPPPP  P PPP PPT T P   PPP P PPPPPP PPPPP  P PP P  PP P   P  P PPTP PP PPPPPPPP  P PPPP   PPPPPPPPPPPP  PPPPPPPPP PPP PTTPPTP PPPPPPPP P                              PP PP  PPPP  PPPPPPPPTPP PPP P   P  PP PP PPPPP  PPP PPPP    P            T                 PPPPPPPPPPPTPPPPPP  PP  PPPPPP PPPPT  PPPP PPPP PPPPP  PP PT PPPP  PPP  PP PPPPP T   PP  PT P  PPPPPPP PPPP  PP PPPP PPPPP       TT   TTT  T            PPPP PPPP   PPPPPPPP  PP PTP PP  PPP      PPPPPP   P PP PPP                                                               TPP  P  PPT PPP PPPPP PPPPPPPPPP PPPP P P PPPPPPPPPPPT  PPPPPP TP PPP  PPP  P   P   PPPPP  PPPPPPP PPPPPPPPPPPPPPPPPPT PPP PPPPPPP PP PP  PPPPP PTPPPP PPPPP  P  PPP PPPPPPPPPP  PPPP     PPPPPP    PP  PP PPPPPPT   PP  PPPPPP  TPP PPPPPPPP P PP PPP PPPPPPP PPP  PPPPPPPP    TP  PPPPPP  PPPP   P PP PP P   PPP T PPP P PPPPPPPPP PT PPP  PPPPPPPPP  PP PPPPPPPTP P PPP  PPPP PP   P P  P PPPP  PT PP P  PPP TPP T  T PPPPP  PPPPPPPPPPPPTPPP PPPPPPPP PP PPPPPPPPPPPP    PPP TPT   P PPPP P  PPPP  P  PP P  PP  PP PPPPPPPPPP TPP     PPPPPPPPPP PPP    P TPPPPPPPP   PP PPPPPPPP PP  PPT T PP  P  PPP T TPP PPP   PP P PPPP PPPP  TP  PPPTPTPT P PP PPPP                  T            PP PPPPPPTTPP    P  PP  PPPPPP  PP  P  PP PPP TPPPPP  T T PPPPPP   PPPP PP   PP  PPP  PPP    PPTPPPPPPPPP         PP PPPPPPP  PPP PP PPPPPP PPPPPP P PP   PPPP PPPP P TPP PP PPT  PPPTP PPPPPPPPP PPPPT PPPPPPPPP  PP PPTP PPTT  P TT PPP   PT  P  PP P  PPPPTTPPP   PPPP PT PPPP  PPPPP  PPPP P  PTP   TPPPT PTPPPPPTT PPPPP PPP     P P PPTT  P PP TP  PPTPPTTPPT   PPPP  T PP   PP P  P  PP   PPTP  PPPPT P T P PPPPP   PPP  PTPPPTPPPPP  PPT  T  PPPPPP  PPP PPPPPPP  P  PPP  PPPP  PP  PPP PP    PPT TPPPPTP TPPPPPPP  PPPPPPPPPPPPP PPP  PP  PPPT    PPTPPPPPPPPT   TP  PPPPPP P PP TPPPPTTTPT                            T TPPPPPPP TPPPPP PP  PPPP PP   P PPP P   PTTP   P PPPP PPPPPP PTPPPPP    P P   PPP PPPTPPP    PPPP" ;
}
