netcdf test_vlen2 {

types:
  int(*) vlen_t;

dimensions:
  d3=3;
  d2=2;
	
variables:
  vlen_t x(d3,d2);  

data:
  x = {1, 3, 5, 7}, {100,200}, {-1,-2},{1, 3, 5, 7}, {100,200}, {-1,-2};
}
