netcdf inttags {
dimensions:
	d = 3 ;
variables:
	byte b(d);
	short s(d);
	int i(d);
data:

 b = -127B, 127b, 255b ;

 s = 32767S, -32766s, 65535s;

 i = -2147483646L, 2147483647l, 4294967295l;
}
