netcdf ref_tst_nul4 {
dimensions:
	n = 8 ;
variables:
	char cdata(n) ;
data:

cdata = "abc\000def" ;
}
