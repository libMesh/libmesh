netcdf test_vlen8 {

types:
  int(*) v_t;

dimensions:
  d1=2;
  d2=2;

variables:
  v_t v1(d1,d2);  

data:

  v1 =
   {1,3,5,7}, {17,19},
   {11,33,55,77}, {717,919};
}

