netcdf inttags4 {
dimensions:
	d = 3 ;
variables:
	ubyte ub(d) ;
	ushort us(d) ;
	uint ui(d) ;
	int64 i64(d) ;
	uint64 ui64(d) ;

// global attributes:
		:attrll = -23232244LL, 1214124123423LL, -2353424234LL ;
data:

 ub = 255, 255, 255 ;

 us = 65534, 65534, 65534 ;

 ui = 4294967294, 4294967294, 4294967294 ;

 i64 = 9223372036854775807, 9223372036854775807, 9223372036854775807 ;

 ui64 = 18446744073709551615, 18446744073709551615, 18446744073709551615 ;
}
