netcdf test {
dimensions:
	\1dim = 1 ;
	dim-name-dashes = 2 ;
	dim.name.dots = 3 ;
	dim+name+plusses = 4 ;
	dim@name@ats = 5 ;
variables:
	float \1var(\1dim) ;
		\1var:\234att = 3 ;
		\1var:att-name-dashes = 4 ;
		\1var:att.name.dots = 5 ;
		\1var:att+name+plusses = 6 ;
		\1var:att@name@ats = 7 ;
	double var-name-dashes ;
	double var.name.dots ;
	double var+name+plusses ;
	double var@name@ats ;

// global attributes:
		:\5Gatt = -1 ;
		:Gatt-name-dashes = -1 ;
		:Gatt.name.dots = -2 ;
		:Gatt+name+plusses = -3 ;
		:Gatt@name@ats = -4 ;
data:

 \1var = _ ;

 var-name-dashes = _ ;

 var.name.dots = _ ;

 var+name+plusses = _ ;

 var@name@ats = _ ;

group: \1g- {
  dimensions:
  	dim\ 1 = 1 ;
  variables:
  	float var\ 1(dim\ 1) ;
  		var\ 1:units\ mks = "km/hour" ;

  // group attributes:
  		:title = "in first group" ;
  data:

   var\ 1 = _ ;
  } // group \1g-
}
