netcdf test_365_day_1900 {
dimensions:
	time = 2300 ;
variables:
	int time(time) ;
		time:units = "days since 1900-1-1" ;
		time:calendar = "365_day" ;
data:

 time = "1900-01-01", "1900-01-02", "1900-01-03", "1900-01-04", "1900-01-05", 
    "1900-01-06", "1900-01-07", "1900-01-08", "1900-01-09", "1900-01-10", 
    "1900-01-11", "1900-01-12", "1900-01-13", "1900-01-14", "1900-01-15", 
    "1900-01-16", "1900-01-17", "1900-01-18", "1900-01-19", "1900-01-20", 
    "1900-01-21", "1900-01-22", "1900-01-23", "1900-01-24", "1900-01-25", 
    "1900-01-26", "1900-01-27", "1900-01-28", "1900-01-29", "1900-01-30", 
    "1900-01-31", "1900-02-01", "1900-02-02", "1900-02-03", "1900-02-04", 
    "1900-02-05", "1900-02-06", "1900-02-07", "1900-02-08", "1900-02-09", 
    "1900-02-10", "1900-02-11", "1900-02-12", "1900-02-13", "1900-02-14", 
    "1900-02-15", "1900-02-16", "1900-02-17", "1900-02-18", "1900-02-19", 
    "1900-02-20", "1900-02-21", "1900-02-22", "1900-02-23", "1900-02-24", 
    "1900-02-25", "1900-02-26", "1900-02-27", "1900-02-28", "1900-03-01", 
    "1900-03-02", "1900-03-03", "1900-03-04", "1900-03-05", "1900-03-06", 
    "1900-03-07", "1900-03-08", "1900-03-09", "1900-03-10", "1900-03-11", 
    "1900-03-12", "1900-03-13", "1900-03-14", "1900-03-15", "1900-03-16", 
    "1900-03-17", "1900-03-18", "1900-03-19", "1900-03-20", "1900-03-21", 
    "1900-03-22", "1900-03-23", "1900-03-24", "1900-03-25", "1900-03-26", 
    "1900-03-27", "1900-03-28", "1900-03-29", "1900-03-30", "1900-03-31", 
    "1900-04-01", "1900-04-02", "1900-04-03", "1900-04-04", "1900-04-05", 
    "1900-04-06", "1900-04-07", "1900-04-08", "1900-04-09", "1900-04-10", 
    "1900-04-11", "1900-04-12", "1900-04-13", "1900-04-14", "1900-04-15", 
    "1900-04-16", "1900-04-17", "1900-04-18", "1900-04-19", "1900-04-20", 
    "1900-04-21", "1900-04-22", "1900-04-23", "1900-04-24", "1900-04-25", 
    "1900-04-26", "1900-04-27", "1900-04-28", "1900-04-29", "1900-04-30", 
    "1900-05-01", "1900-05-02", "1900-05-03", "1900-05-04", "1900-05-05", 
    "1900-05-06", "1900-05-07", "1900-05-08", "1900-05-09", "1900-05-10", 
    "1900-05-11", "1900-05-12", "1900-05-13", "1900-05-14", "1900-05-15", 
    "1900-05-16", "1900-05-17", "1900-05-18", "1900-05-19", "1900-05-20", 
    "1900-05-21", "1900-05-22", "1900-05-23", "1900-05-24", "1900-05-25", 
    "1900-05-26", "1900-05-27", "1900-05-28", "1900-05-29", "1900-05-30", 
    "1900-05-31", "1900-06-01", "1900-06-02", "1900-06-03", "1900-06-04", 
    "1900-06-05", "1900-06-06", "1900-06-07", "1900-06-08", "1900-06-09", 
    "1900-06-10", "1900-06-11", "1900-06-12", "1900-06-13", "1900-06-14", 
    "1900-06-15", "1900-06-16", "1900-06-17", "1900-06-18", "1900-06-19", 
    "1900-06-20", "1900-06-21", "1900-06-22", "1900-06-23", "1900-06-24", 
    "1900-06-25", "1900-06-26", "1900-06-27", "1900-06-28", "1900-06-29", 
    "1900-06-30", "1900-07-01", "1900-07-02", "1900-07-03", "1900-07-04", 
    "1900-07-05", "1900-07-06", "1900-07-07", "1900-07-08", "1900-07-09", 
    "1900-07-10", "1900-07-11", "1900-07-12", "1900-07-13", "1900-07-14", 
    "1900-07-15", "1900-07-16", "1900-07-17", "1900-07-18", "1900-07-19", 
    "1900-07-20", "1900-07-21", "1900-07-22", "1900-07-23", "1900-07-24", 
    "1900-07-25", "1900-07-26", "1900-07-27", "1900-07-28", "1900-07-29", 
    "1900-07-30", "1900-07-31", "1900-08-01", "1900-08-02", "1900-08-03", 
    "1900-08-04", "1900-08-05", "1900-08-06", "1900-08-07", "1900-08-08", 
    "1900-08-09", "1900-08-10", "1900-08-11", "1900-08-12", "1900-08-13", 
    "1900-08-14", "1900-08-15", "1900-08-16", "1900-08-17", "1900-08-18", 
    "1900-08-19", "1900-08-20", "1900-08-21", "1900-08-22", "1900-08-23", 
    "1900-08-24", "1900-08-25", "1900-08-26", "1900-08-27", "1900-08-28", 
    "1900-08-29", "1900-08-30", "1900-08-31", "1900-09-01", "1900-09-02", 
    "1900-09-03", "1900-09-04", "1900-09-05", "1900-09-06", "1900-09-07", 
    "1900-09-08", "1900-09-09", "1900-09-10", "1900-09-11", "1900-09-12", 
    "1900-09-13", "1900-09-14", "1900-09-15", "1900-09-16", "1900-09-17", 
    "1900-09-18", "1900-09-19", "1900-09-20", "1900-09-21", "1900-09-22", 
    "1900-09-23", "1900-09-24", "1900-09-25", "1900-09-26", "1900-09-27", 
    "1900-09-28", "1900-09-29", "1900-09-30", "1900-10-01", "1900-10-02", 
    "1900-10-03", "1900-10-04", "1900-10-05", "1900-10-06", "1900-10-07", 
    "1900-10-08", "1900-10-09", "1900-10-10", "1900-10-11", "1900-10-12", 
    "1900-10-13", "1900-10-14", "1900-10-15", "1900-10-16", "1900-10-17", 
    "1900-10-18", "1900-10-19", "1900-10-20", "1900-10-21", "1900-10-22", 
    "1900-10-23", "1900-10-24", "1900-10-25", "1900-10-26", "1900-10-27", 
    "1900-10-28", "1900-10-29", "1900-10-30", "1900-10-31", "1900-11-01", 
    "1900-11-02", "1900-11-03", "1900-11-04", "1900-11-05", "1900-11-06", 
    "1900-11-07", "1900-11-08", "1900-11-09", "1900-11-10", "1900-11-11", 
    "1900-11-12", "1900-11-13", "1900-11-14", "1900-11-15", "1900-11-16", 
    "1900-11-17", "1900-11-18", "1900-11-19", "1900-11-20", "1900-11-21", 
    "1900-11-22", "1900-11-23", "1900-11-24", "1900-11-25", "1900-11-26", 
    "1900-11-27", "1900-11-28", "1900-11-29", "1900-11-30", "1900-12-01", 
    "1900-12-02", "1900-12-03", "1900-12-04", "1900-12-05", "1900-12-06", 
    "1900-12-07", "1900-12-08", "1900-12-09", "1900-12-10", "1900-12-11", 
    "1900-12-12", "1900-12-13", "1900-12-14", "1900-12-15", "1900-12-16", 
    "1900-12-17", "1900-12-18", "1900-12-19", "1900-12-20", "1900-12-21", 
    "1900-12-22", "1900-12-23", "1900-12-24", "1900-12-25", "1900-12-26", 
    "1900-12-27", "1900-12-28", "1900-12-29", "1900-12-30", "1900-12-31", 
    "1901-01-01", "1901-01-02", "1901-01-03", "1901-01-04", "1901-01-05", 
    "1901-01-06", "1901-01-07", "1901-01-08", "1901-01-09", "1901-01-10", 
    "1901-01-11", "1901-01-12", "1901-01-13", "1901-01-14", "1901-01-15", 
    "1901-01-16", "1901-01-17", "1901-01-18", "1901-01-19", "1901-01-20", 
    "1901-01-21", "1901-01-22", "1901-01-23", "1901-01-24", "1901-01-25", 
    "1901-01-26", "1901-01-27", "1901-01-28", "1901-01-29", "1901-01-30", 
    "1901-01-31", "1901-02-01", "1901-02-02", "1901-02-03", "1901-02-04", 
    "1901-02-05", "1901-02-06", "1901-02-07", "1901-02-08", "1901-02-09", 
    "1901-02-10", "1901-02-11", "1901-02-12", "1901-02-13", "1901-02-14", 
    "1901-02-15", "1901-02-16", "1901-02-17", "1901-02-18", "1901-02-19", 
    "1901-02-20", "1901-02-21", "1901-02-22", "1901-02-23", "1901-02-24", 
    "1901-02-25", "1901-02-26", "1901-02-27", "1901-02-28", "1901-03-01", 
    "1901-03-02", "1901-03-03", "1901-03-04", "1901-03-05", "1901-03-06", 
    "1901-03-07", "1901-03-08", "1901-03-09", "1901-03-10", "1901-03-11", 
    "1901-03-12", "1901-03-13", "1901-03-14", "1901-03-15", "1901-03-16", 
    "1901-03-17", "1901-03-18", "1901-03-19", "1901-03-20", "1901-03-21", 
    "1901-03-22", "1901-03-23", "1901-03-24", "1901-03-25", "1901-03-26", 
    "1901-03-27", "1901-03-28", "1901-03-29", "1901-03-30", "1901-03-31", 
    "1901-04-01", "1901-04-02", "1901-04-03", "1901-04-04", "1901-04-05", 
    "1901-04-06", "1901-04-07", "1901-04-08", "1901-04-09", "1901-04-10", 
    "1901-04-11", "1901-04-12", "1901-04-13", "1901-04-14", "1901-04-15", 
    "1901-04-16", "1901-04-17", "1901-04-18", "1901-04-19", "1901-04-20", 
    "1901-04-21", "1901-04-22", "1901-04-23", "1901-04-24", "1901-04-25", 
    "1901-04-26", "1901-04-27", "1901-04-28", "1901-04-29", "1901-04-30", 
    "1901-05-01", "1901-05-02", "1901-05-03", "1901-05-04", "1901-05-05", 
    "1901-05-06", "1901-05-07", "1901-05-08", "1901-05-09", "1901-05-10", 
    "1901-05-11", "1901-05-12", "1901-05-13", "1901-05-14", "1901-05-15", 
    "1901-05-16", "1901-05-17", "1901-05-18", "1901-05-19", "1901-05-20", 
    "1901-05-21", "1901-05-22", "1901-05-23", "1901-05-24", "1901-05-25", 
    "1901-05-26", "1901-05-27", "1901-05-28", "1901-05-29", "1901-05-30", 
    "1901-05-31", "1901-06-01", "1901-06-02", "1901-06-03", "1901-06-04", 
    "1901-06-05", "1901-06-06", "1901-06-07", "1901-06-08", "1901-06-09", 
    "1901-06-10", "1901-06-11", "1901-06-12", "1901-06-13", "1901-06-14", 
    "1901-06-15", "1901-06-16", "1901-06-17", "1901-06-18", "1901-06-19", 
    "1901-06-20", "1901-06-21", "1901-06-22", "1901-06-23", "1901-06-24", 
    "1901-06-25", "1901-06-26", "1901-06-27", "1901-06-28", "1901-06-29", 
    "1901-06-30", "1901-07-01", "1901-07-02", "1901-07-03", "1901-07-04", 
    "1901-07-05", "1901-07-06", "1901-07-07", "1901-07-08", "1901-07-09", 
    "1901-07-10", "1901-07-11", "1901-07-12", "1901-07-13", "1901-07-14", 
    "1901-07-15", "1901-07-16", "1901-07-17", "1901-07-18", "1901-07-19", 
    "1901-07-20", "1901-07-21", "1901-07-22", "1901-07-23", "1901-07-24", 
    "1901-07-25", "1901-07-26", "1901-07-27", "1901-07-28", "1901-07-29", 
    "1901-07-30", "1901-07-31", "1901-08-01", "1901-08-02", "1901-08-03", 
    "1901-08-04", "1901-08-05", "1901-08-06", "1901-08-07", "1901-08-08", 
    "1901-08-09", "1901-08-10", "1901-08-11", "1901-08-12", "1901-08-13", 
    "1901-08-14", "1901-08-15", "1901-08-16", "1901-08-17", "1901-08-18", 
    "1901-08-19", "1901-08-20", "1901-08-21", "1901-08-22", "1901-08-23", 
    "1901-08-24", "1901-08-25", "1901-08-26", "1901-08-27", "1901-08-28", 
    "1901-08-29", "1901-08-30", "1901-08-31", "1901-09-01", "1901-09-02", 
    "1901-09-03", "1901-09-04", "1901-09-05", "1901-09-06", "1901-09-07", 
    "1901-09-08", "1901-09-09", "1901-09-10", "1901-09-11", "1901-09-12", 
    "1901-09-13", "1901-09-14", "1901-09-15", "1901-09-16", "1901-09-17", 
    "1901-09-18", "1901-09-19", "1901-09-20", "1901-09-21", "1901-09-22", 
    "1901-09-23", "1901-09-24", "1901-09-25", "1901-09-26", "1901-09-27", 
    "1901-09-28", "1901-09-29", "1901-09-30", "1901-10-01", "1901-10-02", 
    "1901-10-03", "1901-10-04", "1901-10-05", "1901-10-06", "1901-10-07", 
    "1901-10-08", "1901-10-09", "1901-10-10", "1901-10-11", "1901-10-12", 
    "1901-10-13", "1901-10-14", "1901-10-15", "1901-10-16", "1901-10-17", 
    "1901-10-18", "1901-10-19", "1901-10-20", "1901-10-21", "1901-10-22", 
    "1901-10-23", "1901-10-24", "1901-10-25", "1901-10-26", "1901-10-27", 
    "1901-10-28", "1901-10-29", "1901-10-30", "1901-10-31", "1901-11-01", 
    "1901-11-02", "1901-11-03", "1901-11-04", "1901-11-05", "1901-11-06", 
    "1901-11-07", "1901-11-08", "1901-11-09", "1901-11-10", "1901-11-11", 
    "1901-11-12", "1901-11-13", "1901-11-14", "1901-11-15", "1901-11-16", 
    "1901-11-17", "1901-11-18", "1901-11-19", "1901-11-20", "1901-11-21", 
    "1901-11-22", "1901-11-23", "1901-11-24", "1901-11-25", "1901-11-26", 
    "1901-11-27", "1901-11-28", "1901-11-29", "1901-11-30", "1901-12-01", 
    "1901-12-02", "1901-12-03", "1901-12-04", "1901-12-05", "1901-12-06", 
    "1901-12-07", "1901-12-08", "1901-12-09", "1901-12-10", "1901-12-11", 
    "1901-12-12", "1901-12-13", "1901-12-14", "1901-12-15", "1901-12-16", 
    "1901-12-17", "1901-12-18", "1901-12-19", "1901-12-20", "1901-12-21", 
    "1901-12-22", "1901-12-23", "1901-12-24", "1901-12-25", "1901-12-26", 
    "1901-12-27", "1901-12-28", "1901-12-29", "1901-12-30", "1901-12-31", 
    "1902-01-01", "1902-01-02", "1902-01-03", "1902-01-04", "1902-01-05", 
    "1902-01-06", "1902-01-07", "1902-01-08", "1902-01-09", "1902-01-10", 
    "1902-01-11", "1902-01-12", "1902-01-13", "1902-01-14", "1902-01-15", 
    "1902-01-16", "1902-01-17", "1902-01-18", "1902-01-19", "1902-01-20", 
    "1902-01-21", "1902-01-22", "1902-01-23", "1902-01-24", "1902-01-25", 
    "1902-01-26", "1902-01-27", "1902-01-28", "1902-01-29", "1902-01-30", 
    "1902-01-31", "1902-02-01", "1902-02-02", "1902-02-03", "1902-02-04", 
    "1902-02-05", "1902-02-06", "1902-02-07", "1902-02-08", "1902-02-09", 
    "1902-02-10", "1902-02-11", "1902-02-12", "1902-02-13", "1902-02-14", 
    "1902-02-15", "1902-02-16", "1902-02-17", "1902-02-18", "1902-02-19", 
    "1902-02-20", "1902-02-21", "1902-02-22", "1902-02-23", "1902-02-24", 
    "1902-02-25", "1902-02-26", "1902-02-27", "1902-02-28", "1902-03-01", 
    "1902-03-02", "1902-03-03", "1902-03-04", "1902-03-05", "1902-03-06", 
    "1902-03-07", "1902-03-08", "1902-03-09", "1902-03-10", "1902-03-11", 
    "1902-03-12", "1902-03-13", "1902-03-14", "1902-03-15", "1902-03-16", 
    "1902-03-17", "1902-03-18", "1902-03-19", "1902-03-20", "1902-03-21", 
    "1902-03-22", "1902-03-23", "1902-03-24", "1902-03-25", "1902-03-26", 
    "1902-03-27", "1902-03-28", "1902-03-29", "1902-03-30", "1902-03-31", 
    "1902-04-01", "1902-04-02", "1902-04-03", "1902-04-04", "1902-04-05", 
    "1902-04-06", "1902-04-07", "1902-04-08", "1902-04-09", "1902-04-10", 
    "1902-04-11", "1902-04-12", "1902-04-13", "1902-04-14", "1902-04-15", 
    "1902-04-16", "1902-04-17", "1902-04-18", "1902-04-19", "1902-04-20", 
    "1902-04-21", "1902-04-22", "1902-04-23", "1902-04-24", "1902-04-25", 
    "1902-04-26", "1902-04-27", "1902-04-28", "1902-04-29", "1902-04-30", 
    "1902-05-01", "1902-05-02", "1902-05-03", "1902-05-04", "1902-05-05", 
    "1902-05-06", "1902-05-07", "1902-05-08", "1902-05-09", "1902-05-10", 
    "1902-05-11", "1902-05-12", "1902-05-13", "1902-05-14", "1902-05-15", 
    "1902-05-16", "1902-05-17", "1902-05-18", "1902-05-19", "1902-05-20", 
    "1902-05-21", "1902-05-22", "1902-05-23", "1902-05-24", "1902-05-25", 
    "1902-05-26", "1902-05-27", "1902-05-28", "1902-05-29", "1902-05-30", 
    "1902-05-31", "1902-06-01", "1902-06-02", "1902-06-03", "1902-06-04", 
    "1902-06-05", "1902-06-06", "1902-06-07", "1902-06-08", "1902-06-09", 
    "1902-06-10", "1902-06-11", "1902-06-12", "1902-06-13", "1902-06-14", 
    "1902-06-15", "1902-06-16", "1902-06-17", "1902-06-18", "1902-06-19", 
    "1902-06-20", "1902-06-21", "1902-06-22", "1902-06-23", "1902-06-24", 
    "1902-06-25", "1902-06-26", "1902-06-27", "1902-06-28", "1902-06-29", 
    "1902-06-30", "1902-07-01", "1902-07-02", "1902-07-03", "1902-07-04", 
    "1902-07-05", "1902-07-06", "1902-07-07", "1902-07-08", "1902-07-09", 
    "1902-07-10", "1902-07-11", "1902-07-12", "1902-07-13", "1902-07-14", 
    "1902-07-15", "1902-07-16", "1902-07-17", "1902-07-18", "1902-07-19", 
    "1902-07-20", "1902-07-21", "1902-07-22", "1902-07-23", "1902-07-24", 
    "1902-07-25", "1902-07-26", "1902-07-27", "1902-07-28", "1902-07-29", 
    "1902-07-30", "1902-07-31", "1902-08-01", "1902-08-02", "1902-08-03", 
    "1902-08-04", "1902-08-05", "1902-08-06", "1902-08-07", "1902-08-08", 
    "1902-08-09", "1902-08-10", "1902-08-11", "1902-08-12", "1902-08-13", 
    "1902-08-14", "1902-08-15", "1902-08-16", "1902-08-17", "1902-08-18", 
    "1902-08-19", "1902-08-20", "1902-08-21", "1902-08-22", "1902-08-23", 
    "1902-08-24", "1902-08-25", "1902-08-26", "1902-08-27", "1902-08-28", 
    "1902-08-29", "1902-08-30", "1902-08-31", "1902-09-01", "1902-09-02", 
    "1902-09-03", "1902-09-04", "1902-09-05", "1902-09-06", "1902-09-07", 
    "1902-09-08", "1902-09-09", "1902-09-10", "1902-09-11", "1902-09-12", 
    "1902-09-13", "1902-09-14", "1902-09-15", "1902-09-16", "1902-09-17", 
    "1902-09-18", "1902-09-19", "1902-09-20", "1902-09-21", "1902-09-22", 
    "1902-09-23", "1902-09-24", "1902-09-25", "1902-09-26", "1902-09-27", 
    "1902-09-28", "1902-09-29", "1902-09-30", "1902-10-01", "1902-10-02", 
    "1902-10-03", "1902-10-04", "1902-10-05", "1902-10-06", "1902-10-07", 
    "1902-10-08", "1902-10-09", "1902-10-10", "1902-10-11", "1902-10-12", 
    "1902-10-13", "1902-10-14", "1902-10-15", "1902-10-16", "1902-10-17", 
    "1902-10-18", "1902-10-19", "1902-10-20", "1902-10-21", "1902-10-22", 
    "1902-10-23", "1902-10-24", "1902-10-25", "1902-10-26", "1902-10-27", 
    "1902-10-28", "1902-10-29", "1902-10-30", "1902-10-31", "1902-11-01", 
    "1902-11-02", "1902-11-03", "1902-11-04", "1902-11-05", "1902-11-06", 
    "1902-11-07", "1902-11-08", "1902-11-09", "1902-11-10", "1902-11-11", 
    "1902-11-12", "1902-11-13", "1902-11-14", "1902-11-15", "1902-11-16", 
    "1902-11-17", "1902-11-18", "1902-11-19", "1902-11-20", "1902-11-21", 
    "1902-11-22", "1902-11-23", "1902-11-24", "1902-11-25", "1902-11-26", 
    "1902-11-27", "1902-11-28", "1902-11-29", "1902-11-30", "1902-12-01", 
    "1902-12-02", "1902-12-03", "1902-12-04", "1902-12-05", "1902-12-06", 
    "1902-12-07", "1902-12-08", "1902-12-09", "1902-12-10", "1902-12-11", 
    "1902-12-12", "1902-12-13", "1902-12-14", "1902-12-15", "1902-12-16", 
    "1902-12-17", "1902-12-18", "1902-12-19", "1902-12-20", "1902-12-21", 
    "1902-12-22", "1902-12-23", "1902-12-24", "1902-12-25", "1902-12-26", 
    "1902-12-27", "1902-12-28", "1902-12-29", "1902-12-30", "1902-12-31", 
    "1903-01-01", "1903-01-02", "1903-01-03", "1903-01-04", "1903-01-05", 
    "1903-01-06", "1903-01-07", "1903-01-08", "1903-01-09", "1903-01-10", 
    "1903-01-11", "1903-01-12", "1903-01-13", "1903-01-14", "1903-01-15", 
    "1903-01-16", "1903-01-17", "1903-01-18", "1903-01-19", "1903-01-20", 
    "1903-01-21", "1903-01-22", "1903-01-23", "1903-01-24", "1903-01-25", 
    "1903-01-26", "1903-01-27", "1903-01-28", "1903-01-29", "1903-01-30", 
    "1903-01-31", "1903-02-01", "1903-02-02", "1903-02-03", "1903-02-04", 
    "1903-02-05", "1903-02-06", "1903-02-07", "1903-02-08", "1903-02-09", 
    "1903-02-10", "1903-02-11", "1903-02-12", "1903-02-13", "1903-02-14", 
    "1903-02-15", "1903-02-16", "1903-02-17", "1903-02-18", "1903-02-19", 
    "1903-02-20", "1903-02-21", "1903-02-22", "1903-02-23", "1903-02-24", 
    "1903-02-25", "1903-02-26", "1903-02-27", "1903-02-28", "1903-03-01", 
    "1903-03-02", "1903-03-03", "1903-03-04", "1903-03-05", "1903-03-06", 
    "1903-03-07", "1903-03-08", "1903-03-09", "1903-03-10", "1903-03-11", 
    "1903-03-12", "1903-03-13", "1903-03-14", "1903-03-15", "1903-03-16", 
    "1903-03-17", "1903-03-18", "1903-03-19", "1903-03-20", "1903-03-21", 
    "1903-03-22", "1903-03-23", "1903-03-24", "1903-03-25", "1903-03-26", 
    "1903-03-27", "1903-03-28", "1903-03-29", "1903-03-30", "1903-03-31", 
    "1903-04-01", "1903-04-02", "1903-04-03", "1903-04-04", "1903-04-05", 
    "1903-04-06", "1903-04-07", "1903-04-08", "1903-04-09", "1903-04-10", 
    "1903-04-11", "1903-04-12", "1903-04-13", "1903-04-14", "1903-04-15", 
    "1903-04-16", "1903-04-17", "1903-04-18", "1903-04-19", "1903-04-20", 
    "1903-04-21", "1903-04-22", "1903-04-23", "1903-04-24", "1903-04-25", 
    "1903-04-26", "1903-04-27", "1903-04-28", "1903-04-29", "1903-04-30", 
    "1903-05-01", "1903-05-02", "1903-05-03", "1903-05-04", "1903-05-05", 
    "1903-05-06", "1903-05-07", "1903-05-08", "1903-05-09", "1903-05-10", 
    "1903-05-11", "1903-05-12", "1903-05-13", "1903-05-14", "1903-05-15", 
    "1903-05-16", "1903-05-17", "1903-05-18", "1903-05-19", "1903-05-20", 
    "1903-05-21", "1903-05-22", "1903-05-23", "1903-05-24", "1903-05-25", 
    "1903-05-26", "1903-05-27", "1903-05-28", "1903-05-29", "1903-05-30", 
    "1903-05-31", "1903-06-01", "1903-06-02", "1903-06-03", "1903-06-04", 
    "1903-06-05", "1903-06-06", "1903-06-07", "1903-06-08", "1903-06-09", 
    "1903-06-10", "1903-06-11", "1903-06-12", "1903-06-13", "1903-06-14", 
    "1903-06-15", "1903-06-16", "1903-06-17", "1903-06-18", "1903-06-19", 
    "1903-06-20", "1903-06-21", "1903-06-22", "1903-06-23", "1903-06-24", 
    "1903-06-25", "1903-06-26", "1903-06-27", "1903-06-28", "1903-06-29", 
    "1903-06-30", "1903-07-01", "1903-07-02", "1903-07-03", "1903-07-04", 
    "1903-07-05", "1903-07-06", "1903-07-07", "1903-07-08", "1903-07-09", 
    "1903-07-10", "1903-07-11", "1903-07-12", "1903-07-13", "1903-07-14", 
    "1903-07-15", "1903-07-16", "1903-07-17", "1903-07-18", "1903-07-19", 
    "1903-07-20", "1903-07-21", "1903-07-22", "1903-07-23", "1903-07-24", 
    "1903-07-25", "1903-07-26", "1903-07-27", "1903-07-28", "1903-07-29", 
    "1903-07-30", "1903-07-31", "1903-08-01", "1903-08-02", "1903-08-03", 
    "1903-08-04", "1903-08-05", "1903-08-06", "1903-08-07", "1903-08-08", 
    "1903-08-09", "1903-08-10", "1903-08-11", "1903-08-12", "1903-08-13", 
    "1903-08-14", "1903-08-15", "1903-08-16", "1903-08-17", "1903-08-18", 
    "1903-08-19", "1903-08-20", "1903-08-21", "1903-08-22", "1903-08-23", 
    "1903-08-24", "1903-08-25", "1903-08-26", "1903-08-27", "1903-08-28", 
    "1903-08-29", "1903-08-30", "1903-08-31", "1903-09-01", "1903-09-02", 
    "1903-09-03", "1903-09-04", "1903-09-05", "1903-09-06", "1903-09-07", 
    "1903-09-08", "1903-09-09", "1903-09-10", "1903-09-11", "1903-09-12", 
    "1903-09-13", "1903-09-14", "1903-09-15", "1903-09-16", "1903-09-17", 
    "1903-09-18", "1903-09-19", "1903-09-20", "1903-09-21", "1903-09-22", 
    "1903-09-23", "1903-09-24", "1903-09-25", "1903-09-26", "1903-09-27", 
    "1903-09-28", "1903-09-29", "1903-09-30", "1903-10-01", "1903-10-02", 
    "1903-10-03", "1903-10-04", "1903-10-05", "1903-10-06", "1903-10-07", 
    "1903-10-08", "1903-10-09", "1903-10-10", "1903-10-11", "1903-10-12", 
    "1903-10-13", "1903-10-14", "1903-10-15", "1903-10-16", "1903-10-17", 
    "1903-10-18", "1903-10-19", "1903-10-20", "1903-10-21", "1903-10-22", 
    "1903-10-23", "1903-10-24", "1903-10-25", "1903-10-26", "1903-10-27", 
    "1903-10-28", "1903-10-29", "1903-10-30", "1903-10-31", "1903-11-01", 
    "1903-11-02", "1903-11-03", "1903-11-04", "1903-11-05", "1903-11-06", 
    "1903-11-07", "1903-11-08", "1903-11-09", "1903-11-10", "1903-11-11", 
    "1903-11-12", "1903-11-13", "1903-11-14", "1903-11-15", "1903-11-16", 
    "1903-11-17", "1903-11-18", "1903-11-19", "1903-11-20", "1903-11-21", 
    "1903-11-22", "1903-11-23", "1903-11-24", "1903-11-25", "1903-11-26", 
    "1903-11-27", "1903-11-28", "1903-11-29", "1903-11-30", "1903-12-01", 
    "1903-12-02", "1903-12-03", "1903-12-04", "1903-12-05", "1903-12-06", 
    "1903-12-07", "1903-12-08", "1903-12-09", "1903-12-10", "1903-12-11", 
    "1903-12-12", "1903-12-13", "1903-12-14", "1903-12-15", "1903-12-16", 
    "1903-12-17", "1903-12-18", "1903-12-19", "1903-12-20", "1903-12-21", 
    "1903-12-22", "1903-12-23", "1903-12-24", "1903-12-25", "1903-12-26", 
    "1903-12-27", "1903-12-28", "1903-12-29", "1903-12-30", "1903-12-31", 
    "1904-01-01", "1904-01-02", "1904-01-03", "1904-01-04", "1904-01-05", 
    "1904-01-06", "1904-01-07", "1904-01-08", "1904-01-09", "1904-01-10", 
    "1904-01-11", "1904-01-12", "1904-01-13", "1904-01-14", "1904-01-15", 
    "1904-01-16", "1904-01-17", "1904-01-18", "1904-01-19", "1904-01-20", 
    "1904-01-21", "1904-01-22", "1904-01-23", "1904-01-24", "1904-01-25", 
    "1904-01-26", "1904-01-27", "1904-01-28", "1904-01-29", "1904-01-30", 
    "1904-01-31", "1904-02-01", "1904-02-02", "1904-02-03", "1904-02-04", 
    "1904-02-05", "1904-02-06", "1904-02-07", "1904-02-08", "1904-02-09", 
    "1904-02-10", "1904-02-11", "1904-02-12", "1904-02-13", "1904-02-14", 
    "1904-02-15", "1904-02-16", "1904-02-17", "1904-02-18", "1904-02-19", 
    "1904-02-20", "1904-02-21", "1904-02-22", "1904-02-23", "1904-02-24", 
    "1904-02-25", "1904-02-26", "1904-02-27", "1904-02-28", "1904-03-01", 
    "1904-03-02", "1904-03-03", "1904-03-04", "1904-03-05", "1904-03-06", 
    "1904-03-07", "1904-03-08", "1904-03-09", "1904-03-10", "1904-03-11", 
    "1904-03-12", "1904-03-13", "1904-03-14", "1904-03-15", "1904-03-16", 
    "1904-03-17", "1904-03-18", "1904-03-19", "1904-03-20", "1904-03-21", 
    "1904-03-22", "1904-03-23", "1904-03-24", "1904-03-25", "1904-03-26", 
    "1904-03-27", "1904-03-28", "1904-03-29", "1904-03-30", "1904-03-31", 
    "1904-04-01", "1904-04-02", "1904-04-03", "1904-04-04", "1904-04-05", 
    "1904-04-06", "1904-04-07", "1904-04-08", "1904-04-09", "1904-04-10", 
    "1904-04-11", "1904-04-12", "1904-04-13", "1904-04-14", "1904-04-15", 
    "1904-04-16", "1904-04-17", "1904-04-18", "1904-04-19", "1904-04-20", 
    "1904-04-21", "1904-04-22", "1904-04-23", "1904-04-24", "1904-04-25", 
    "1904-04-26", "1904-04-27", "1904-04-28", "1904-04-29", "1904-04-30", 
    "1904-05-01", "1904-05-02", "1904-05-03", "1904-05-04", "1904-05-05", 
    "1904-05-06", "1904-05-07", "1904-05-08", "1904-05-09", "1904-05-10", 
    "1904-05-11", "1904-05-12", "1904-05-13", "1904-05-14", "1904-05-15", 
    "1904-05-16", "1904-05-17", "1904-05-18", "1904-05-19", "1904-05-20", 
    "1904-05-21", "1904-05-22", "1904-05-23", "1904-05-24", "1904-05-25", 
    "1904-05-26", "1904-05-27", "1904-05-28", "1904-05-29", "1904-05-30", 
    "1904-05-31", "1904-06-01", "1904-06-02", "1904-06-03", "1904-06-04", 
    "1904-06-05", "1904-06-06", "1904-06-07", "1904-06-08", "1904-06-09", 
    "1904-06-10", "1904-06-11", "1904-06-12", "1904-06-13", "1904-06-14", 
    "1904-06-15", "1904-06-16", "1904-06-17", "1904-06-18", "1904-06-19", 
    "1904-06-20", "1904-06-21", "1904-06-22", "1904-06-23", "1904-06-24", 
    "1904-06-25", "1904-06-26", "1904-06-27", "1904-06-28", "1904-06-29", 
    "1904-06-30", "1904-07-01", "1904-07-02", "1904-07-03", "1904-07-04", 
    "1904-07-05", "1904-07-06", "1904-07-07", "1904-07-08", "1904-07-09", 
    "1904-07-10", "1904-07-11", "1904-07-12", "1904-07-13", "1904-07-14", 
    "1904-07-15", "1904-07-16", "1904-07-17", "1904-07-18", "1904-07-19", 
    "1904-07-20", "1904-07-21", "1904-07-22", "1904-07-23", "1904-07-24", 
    "1904-07-25", "1904-07-26", "1904-07-27", "1904-07-28", "1904-07-29", 
    "1904-07-30", "1904-07-31", "1904-08-01", "1904-08-02", "1904-08-03", 
    "1904-08-04", "1904-08-05", "1904-08-06", "1904-08-07", "1904-08-08", 
    "1904-08-09", "1904-08-10", "1904-08-11", "1904-08-12", "1904-08-13", 
    "1904-08-14", "1904-08-15", "1904-08-16", "1904-08-17", "1904-08-18", 
    "1904-08-19", "1904-08-20", "1904-08-21", "1904-08-22", "1904-08-23", 
    "1904-08-24", "1904-08-25", "1904-08-26", "1904-08-27", "1904-08-28", 
    "1904-08-29", "1904-08-30", "1904-08-31", "1904-09-01", "1904-09-02", 
    "1904-09-03", "1904-09-04", "1904-09-05", "1904-09-06", "1904-09-07", 
    "1904-09-08", "1904-09-09", "1904-09-10", "1904-09-11", "1904-09-12", 
    "1904-09-13", "1904-09-14", "1904-09-15", "1904-09-16", "1904-09-17", 
    "1904-09-18", "1904-09-19", "1904-09-20", "1904-09-21", "1904-09-22", 
    "1904-09-23", "1904-09-24", "1904-09-25", "1904-09-26", "1904-09-27", 
    "1904-09-28", "1904-09-29", "1904-09-30", "1904-10-01", "1904-10-02", 
    "1904-10-03", "1904-10-04", "1904-10-05", "1904-10-06", "1904-10-07", 
    "1904-10-08", "1904-10-09", "1904-10-10", "1904-10-11", "1904-10-12", 
    "1904-10-13", "1904-10-14", "1904-10-15", "1904-10-16", "1904-10-17", 
    "1904-10-18", "1904-10-19", "1904-10-20", "1904-10-21", "1904-10-22", 
    "1904-10-23", "1904-10-24", "1904-10-25", "1904-10-26", "1904-10-27", 
    "1904-10-28", "1904-10-29", "1904-10-30", "1904-10-31", "1904-11-01", 
    "1904-11-02", "1904-11-03", "1904-11-04", "1904-11-05", "1904-11-06", 
    "1904-11-07", "1904-11-08", "1904-11-09", "1904-11-10", "1904-11-11", 
    "1904-11-12", "1904-11-13", "1904-11-14", "1904-11-15", "1904-11-16", 
    "1904-11-17", "1904-11-18", "1904-11-19", "1904-11-20", "1904-11-21", 
    "1904-11-22", "1904-11-23", "1904-11-24", "1904-11-25", "1904-11-26", 
    "1904-11-27", "1904-11-28", "1904-11-29", "1904-11-30", "1904-12-01", 
    "1904-12-02", "1904-12-03", "1904-12-04", "1904-12-05", "1904-12-06", 
    "1904-12-07", "1904-12-08", "1904-12-09", "1904-12-10", "1904-12-11", 
    "1904-12-12", "1904-12-13", "1904-12-14", "1904-12-15", "1904-12-16", 
    "1904-12-17", "1904-12-18", "1904-12-19", "1904-12-20", "1904-12-21", 
    "1904-12-22", "1904-12-23", "1904-12-24", "1904-12-25", "1904-12-26", 
    "1904-12-27", "1904-12-28", "1904-12-29", "1904-12-30", "1904-12-31", 
    "1905-01-01", "1905-01-02", "1905-01-03", "1905-01-04", "1905-01-05", 
    "1905-01-06", "1905-01-07", "1905-01-08", "1905-01-09", "1905-01-10", 
    "1905-01-11", "1905-01-12", "1905-01-13", "1905-01-14", "1905-01-15", 
    "1905-01-16", "1905-01-17", "1905-01-18", "1905-01-19", "1905-01-20", 
    "1905-01-21", "1905-01-22", "1905-01-23", "1905-01-24", "1905-01-25", 
    "1905-01-26", "1905-01-27", "1905-01-28", "1905-01-29", "1905-01-30", 
    "1905-01-31", "1905-02-01", "1905-02-02", "1905-02-03", "1905-02-04", 
    "1905-02-05", "1905-02-06", "1905-02-07", "1905-02-08", "1905-02-09", 
    "1905-02-10", "1905-02-11", "1905-02-12", "1905-02-13", "1905-02-14", 
    "1905-02-15", "1905-02-16", "1905-02-17", "1905-02-18", "1905-02-19", 
    "1905-02-20", "1905-02-21", "1905-02-22", "1905-02-23", "1905-02-24", 
    "1905-02-25", "1905-02-26", "1905-02-27", "1905-02-28", "1905-03-01", 
    "1905-03-02", "1905-03-03", "1905-03-04", "1905-03-05", "1905-03-06", 
    "1905-03-07", "1905-03-08", "1905-03-09", "1905-03-10", "1905-03-11", 
    "1905-03-12", "1905-03-13", "1905-03-14", "1905-03-15", "1905-03-16", 
    "1905-03-17", "1905-03-18", "1905-03-19", "1905-03-20", "1905-03-21", 
    "1905-03-22", "1905-03-23", "1905-03-24", "1905-03-25", "1905-03-26", 
    "1905-03-27", "1905-03-28", "1905-03-29", "1905-03-30", "1905-03-31", 
    "1905-04-01", "1905-04-02", "1905-04-03", "1905-04-04", "1905-04-05", 
    "1905-04-06", "1905-04-07", "1905-04-08", "1905-04-09", "1905-04-10", 
    "1905-04-11", "1905-04-12", "1905-04-13", "1905-04-14", "1905-04-15", 
    "1905-04-16", "1905-04-17", "1905-04-18", "1905-04-19", "1905-04-20", 
    "1905-04-21", "1905-04-22", "1905-04-23", "1905-04-24", "1905-04-25", 
    "1905-04-26", "1905-04-27", "1905-04-28", "1905-04-29", "1905-04-30", 
    "1905-05-01", "1905-05-02", "1905-05-03", "1905-05-04", "1905-05-05", 
    "1905-05-06", "1905-05-07", "1905-05-08", "1905-05-09", "1905-05-10", 
    "1905-05-11", "1905-05-12", "1905-05-13", "1905-05-14", "1905-05-15", 
    "1905-05-16", "1905-05-17", "1905-05-18", "1905-05-19", "1905-05-20", 
    "1905-05-21", "1905-05-22", "1905-05-23", "1905-05-24", "1905-05-25", 
    "1905-05-26", "1905-05-27", "1905-05-28", "1905-05-29", "1905-05-30", 
    "1905-05-31", "1905-06-01", "1905-06-02", "1905-06-03", "1905-06-04", 
    "1905-06-05", "1905-06-06", "1905-06-07", "1905-06-08", "1905-06-09", 
    "1905-06-10", "1905-06-11", "1905-06-12", "1905-06-13", "1905-06-14", 
    "1905-06-15", "1905-06-16", "1905-06-17", "1905-06-18", "1905-06-19", 
    "1905-06-20", "1905-06-21", "1905-06-22", "1905-06-23", "1905-06-24", 
    "1905-06-25", "1905-06-26", "1905-06-27", "1905-06-28", "1905-06-29", 
    "1905-06-30", "1905-07-01", "1905-07-02", "1905-07-03", "1905-07-04", 
    "1905-07-05", "1905-07-06", "1905-07-07", "1905-07-08", "1905-07-09", 
    "1905-07-10", "1905-07-11", "1905-07-12", "1905-07-13", "1905-07-14", 
    "1905-07-15", "1905-07-16", "1905-07-17", "1905-07-18", "1905-07-19", 
    "1905-07-20", "1905-07-21", "1905-07-22", "1905-07-23", "1905-07-24", 
    "1905-07-25", "1905-07-26", "1905-07-27", "1905-07-28", "1905-07-29", 
    "1905-07-30", "1905-07-31", "1905-08-01", "1905-08-02", "1905-08-03", 
    "1905-08-04", "1905-08-05", "1905-08-06", "1905-08-07", "1905-08-08", 
    "1905-08-09", "1905-08-10", "1905-08-11", "1905-08-12", "1905-08-13", 
    "1905-08-14", "1905-08-15", "1905-08-16", "1905-08-17", "1905-08-18", 
    "1905-08-19", "1905-08-20", "1905-08-21", "1905-08-22", "1905-08-23", 
    "1905-08-24", "1905-08-25", "1905-08-26", "1905-08-27", "1905-08-28", 
    "1905-08-29", "1905-08-30", "1905-08-31", "1905-09-01", "1905-09-02", 
    "1905-09-03", "1905-09-04", "1905-09-05", "1905-09-06", "1905-09-07", 
    "1905-09-08", "1905-09-09", "1905-09-10", "1905-09-11", "1905-09-12", 
    "1905-09-13", "1905-09-14", "1905-09-15", "1905-09-16", "1905-09-17", 
    "1905-09-18", "1905-09-19", "1905-09-20", "1905-09-21", "1905-09-22", 
    "1905-09-23", "1905-09-24", "1905-09-25", "1905-09-26", "1905-09-27", 
    "1905-09-28", "1905-09-29", "1905-09-30", "1905-10-01", "1905-10-02", 
    "1905-10-03", "1905-10-04", "1905-10-05", "1905-10-06", "1905-10-07", 
    "1905-10-08", "1905-10-09", "1905-10-10", "1905-10-11", "1905-10-12", 
    "1905-10-13", "1905-10-14", "1905-10-15", "1905-10-16", "1905-10-17", 
    "1905-10-18", "1905-10-19", "1905-10-20", "1905-10-21", "1905-10-22", 
    "1905-10-23", "1905-10-24", "1905-10-25", "1905-10-26", "1905-10-27", 
    "1905-10-28", "1905-10-29", "1905-10-30", "1905-10-31", "1905-11-01", 
    "1905-11-02", "1905-11-03", "1905-11-04", "1905-11-05", "1905-11-06", 
    "1905-11-07", "1905-11-08", "1905-11-09", "1905-11-10", "1905-11-11", 
    "1905-11-12", "1905-11-13", "1905-11-14", "1905-11-15", "1905-11-16", 
    "1905-11-17", "1905-11-18", "1905-11-19", "1905-11-20", "1905-11-21", 
    "1905-11-22", "1905-11-23", "1905-11-24", "1905-11-25", "1905-11-26", 
    "1905-11-27", "1905-11-28", "1905-11-29", "1905-11-30", "1905-12-01", 
    "1905-12-02", "1905-12-03", "1905-12-04", "1905-12-05", "1905-12-06", 
    "1905-12-07", "1905-12-08", "1905-12-09", "1905-12-10", "1905-12-11", 
    "1905-12-12", "1905-12-13", "1905-12-14", "1905-12-15", "1905-12-16", 
    "1905-12-17", "1905-12-18", "1905-12-19", "1905-12-20", "1905-12-21", 
    "1905-12-22", "1905-12-23", "1905-12-24", "1905-12-25", "1905-12-26", 
    "1905-12-27", "1905-12-28", "1905-12-29", "1905-12-30", "1905-12-31", 
    "1906-01-01", "1906-01-02", "1906-01-03", "1906-01-04", "1906-01-05", 
    "1906-01-06", "1906-01-07", "1906-01-08", "1906-01-09", "1906-01-10", 
    "1906-01-11", "1906-01-12", "1906-01-13", "1906-01-14", "1906-01-15", 
    "1906-01-16", "1906-01-17", "1906-01-18", "1906-01-19", "1906-01-20", 
    "1906-01-21", "1906-01-22", "1906-01-23", "1906-01-24", "1906-01-25", 
    "1906-01-26", "1906-01-27", "1906-01-28", "1906-01-29", "1906-01-30", 
    "1906-01-31", "1906-02-01", "1906-02-02", "1906-02-03", "1906-02-04", 
    "1906-02-05", "1906-02-06", "1906-02-07", "1906-02-08", "1906-02-09", 
    "1906-02-10", "1906-02-11", "1906-02-12", "1906-02-13", "1906-02-14", 
    "1906-02-15", "1906-02-16", "1906-02-17", "1906-02-18", "1906-02-19", 
    "1906-02-20", "1906-02-21", "1906-02-22", "1906-02-23", "1906-02-24", 
    "1906-02-25", "1906-02-26", "1906-02-27", "1906-02-28", "1906-03-01", 
    "1906-03-02", "1906-03-03", "1906-03-04", "1906-03-05", "1906-03-06", 
    "1906-03-07", "1906-03-08", "1906-03-09", "1906-03-10", "1906-03-11", 
    "1906-03-12", "1906-03-13", "1906-03-14", "1906-03-15", "1906-03-16", 
    "1906-03-17", "1906-03-18", "1906-03-19", "1906-03-20", "1906-03-21", 
    "1906-03-22", "1906-03-23", "1906-03-24", "1906-03-25", "1906-03-26", 
    "1906-03-27", "1906-03-28", "1906-03-29", "1906-03-30", "1906-03-31", 
    "1906-04-01", "1906-04-02", "1906-04-03", "1906-04-04", "1906-04-05", 
    "1906-04-06", "1906-04-07", "1906-04-08", "1906-04-09", "1906-04-10", 
    "1906-04-11", "1906-04-12", "1906-04-13", "1906-04-14", "1906-04-15", 
    "1906-04-16", "1906-04-17", "1906-04-18", "1906-04-19", "1906-04-20" ;
}
