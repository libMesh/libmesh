netcdf test_struct_array {
types:
    compound c_t {
      int x ;
      int y ;
    }; // c_t
dimensions:
 dx = 4;
 dy = 3;
variables:
  c_t s(dx,dy);
data:
 s =
/*[0][0..2]*/  {1, -1}, {17, 37}, {-32767, 32767},
/*[1][0..2]*/  {-1, 3}, {-2, 2}, {-3, 1},
/*[2][0..2]*/  {-4, 12}, {-8, 8}, {-12, 4},
/*[3][0..2]*/  {-5, 15}, {-10, 10}, {-15, 5} ;
}
